`default_nettype none

module fsqrt
    ( input wire [31:0] x,
      output wire [31:0] y,
      input wire clk,
      input wire rstn
);
    wire en;
    wire we;
    wire rst;
    wire [35:0] din;

    assign en = 1;
    assign we = 0;
    assign rst = 0;
    assign din = 0;

    wire s;
    wire [7:0] e;
    wire [22:0] m;
    wire [35:0] val;
    wire [9:0] key;

    wire [22:0] c;
    wire [29:0] cor_n;

    reg s_reg;
    reg s_reg2;
    reg [7:0] e_reg;
    reg [7:0] e_reg2;
    reg [22:0] m_reg;
    reg [29:0] cor_n_reg;
    reg [22:0] c_reg;
    reg [9:0] key_reg;
    reg [35:0] val_reg;

    assign s = x[31];
    assign e = x[30:23];
    assign m = x[22:0];
    assign key = x[23:14];

    fsqrt_table u1(clk, en, we, rst, key, din, val);
    fsqrt_1st u2(m_reg, key_reg, val, c, cor_n);
    fsqrt_2nd u3(s_reg2, e_reg2, c_reg, cor_n_reg, y);

    always @(posedge clk) begin
        s_reg <= s;
        s_reg2 <= s_reg;
        e_reg <= e;
        e_reg2 <= e_reg;
        m_reg <= m;
        key_reg <= key;
        val_reg <= val;
        c_reg <= c;
        cor_n_reg <= cor_n;
    end

endmodule


module fsqrt_1st
    (input wire [22:0] m,
     input wire [9:0] key,
     input wire [35:0] val,
     output wire [22:0] c,
     output wire [29:0] cor_n);

    wire [13:0] d;
    wire [13:0] a1;
    wire [14:0] a2;

    assign c = val[35:13];
    assign d = {1'b1, val[12:0]};
    assign a1 = m[13:0];
    assign a2 = a1 << 1;
    assign cor_n = (key < 10'd512) ? a2 * d : a1 * d;

endmodule

module fsqrt_2nd
    (input wire s,
     input wire [7:0] e,
     input wire [22:0] c,
     input wire [29:0] cor_n,
     output wire [31:0] y);

    wire [22:0] ans_m;
    wire [22:0] m1;
    wire [8:0] e0;
    wire [7:0] ans_e;
    wire [14:0] cor;

    assign cor = cor_n >> 15;
    assign e0 = e + 8'd127;
    assign ans_e = e0[8:1];
    assign m1 = c + cor;
    assign ans_m = (e == 0) ? 0 : m1;
    assign y = (e == 0) ? {s, 8'b0, ans_m} : {s, ans_e, ans_m};

endmodule



module fsqrt_table
(
    input wire clk,
    input wire en,
    input wire we,
    input wire rst,
    input wire [9:0] addr,
    input wire [35:0] di,
    output reg [35:0] dout
);

    reg [35:0] fsqrt_table [1023:0];

initial
    begin
        fsqrt_table[1023] = 36'h69DCA2D45;
        fsqrt_table[1022] = 36'h69AF58D4B;
        fsqrt_table[1021] = 36'h69820AD4E;
        fsqrt_table[1020] = 36'h6954B4D55;
        fsqrt_table[1019] = 36'h69275AD5A;
        fsqrt_table[1018] = 36'h68F9FAD5F;
        fsqrt_table[1017] = 36'h68CC94D64;
        fsqrt_table[1016] = 36'h689F28D6A;
        fsqrt_table[1015] = 36'h6871B6D70;
        fsqrt_table[1014] = 36'h68443ED77;
        fsqrt_table[1013] = 36'h6816C2D7B;
        fsqrt_table[1012] = 36'h67E93ED83;
        fsqrt_table[1011] = 36'h67BBB6D87;
        fsqrt_table[1010] = 36'h678E28D8D;
        fsqrt_table[1009] = 36'h676094D92;
        fsqrt_table[1008] = 36'h6732FAD98;
        fsqrt_table[1007] = 36'h67055AD9E;
        fsqrt_table[1006] = 36'h66D7B4DA5;
        fsqrt_table[1005] = 36'h66AA08DAC;
        fsqrt_table[1004] = 36'h667C58DB0;
        fsqrt_table[1003] = 36'h664EA0DB7;
        fsqrt_table[1002] = 36'h6620E4DBC;
        fsqrt_table[1001] = 36'h65F320DC4;
        fsqrt_table[1000] = 36'h65C558DC9;
        fsqrt_table[999] = 36'h65978ADCE;
        fsqrt_table[998] = 36'h6569B6DD4;
        fsqrt_table[997] = 36'h653BDCDD9;
        fsqrt_table[996] = 36'h650DFCDDF;
        fsqrt_table[995] = 36'h64E016DE5;
        fsqrt_table[994] = 36'h64B22ADEB;
        fsqrt_table[993] = 36'h648438DF2;
        fsqrt_table[992] = 36'h645640DF8;
        fsqrt_table[991] = 36'h642842DFF;
        fsqrt_table[990] = 36'h63FA40E02;
        fsqrt_table[989] = 36'h63CC36E09;
        fsqrt_table[988] = 36'h639E26E10;
        fsqrt_table[987] = 36'h637012E14;
        fsqrt_table[986] = 36'h6341F6E1B;
        fsqrt_table[985] = 36'h6313D4E22;
        fsqrt_table[984] = 36'h62E5ACE29;
        fsqrt_table[983] = 36'h62B780E2D;
        fsqrt_table[982] = 36'h62894CE34;
        fsqrt_table[981] = 36'h625B12E3B;
        fsqrt_table[980] = 36'h622CD4E3E;
        fsqrt_table[979] = 36'h61FE8EE45;
        fsqrt_table[978] = 36'h61D042E4C;
        fsqrt_table[977] = 36'h61A1F0E53;
        fsqrt_table[976] = 36'h61739AE56;
        fsqrt_table[975] = 36'h61453CE5D;
        fsqrt_table[974] = 36'h6116D8E63;
        fsqrt_table[973] = 36'h60E86EE69;
        fsqrt_table[972] = 36'h60B9FEE6F;
        fsqrt_table[971] = 36'h608B88E75;
        fsqrt_table[970] = 36'h605D0CE7B;
        fsqrt_table[969] = 36'h602E8AE81;
        fsqrt_table[968] = 36'h600000E89;
        fsqrt_table[967] = 36'h5FD172E8E;
        fsqrt_table[966] = 36'h5FA2DCE96;
        fsqrt_table[965] = 36'h5F7442E9A;
        fsqrt_table[964] = 36'h5F45A0EA2;
        fsqrt_table[963] = 36'h5F16F8EA9;
        fsqrt_table[962] = 36'h5EE84CEAC;
        fsqrt_table[961] = 36'h5EB998EB3;
        fsqrt_table[960] = 36'h5E8ADEEB9;
        fsqrt_table[959] = 36'h5E5C1CEC2;
        fsqrt_table[958] = 36'h5E2D56EC7;
        fsqrt_table[957] = 36'h5DFE8AECC;
        fsqrt_table[956] = 36'h5DCFB6ED4;
        fsqrt_table[955] = 36'h5DA0DEED8;
        fsqrt_table[954] = 36'h5D71FEEDF;
        fsqrt_table[953] = 36'h5D4318EE5;
        fsqrt_table[952] = 36'h5D142CEEB;
        fsqrt_table[951] = 36'h5CE53AEF1;
        fsqrt_table[950] = 36'h5CB640EF9;
        fsqrt_table[949] = 36'h5C8742EFE;
        fsqrt_table[948] = 36'h5C583CF05;
        fsqrt_table[947] = 36'h5C2930F0B;
        fsqrt_table[946] = 36'h5BFA1EF11;
        fsqrt_table[945] = 36'h5BCB06F17;
        fsqrt_table[944] = 36'h5B9BE6F1F;
        fsqrt_table[943] = 36'h5B6CC0F26;
        fsqrt_table[942] = 36'h5B3D96F2A;
        fsqrt_table[941] = 36'h5B0E62F33;
        fsqrt_table[940] = 36'h5ADF2AF39;
        fsqrt_table[939] = 36'h5AAFECF3E;
        fsqrt_table[938] = 36'h5A80A6F45;
        fsqrt_table[937] = 36'h5A515AF4B;
        fsqrt_table[936] = 36'h5A2208F51;
        fsqrt_table[935] = 36'h59F2AEF5A;
        fsqrt_table[934] = 36'h59C350F5E;
        fsqrt_table[933] = 36'h5993EAF65;
        fsqrt_table[932] = 36'h59647EF6B;
        fsqrt_table[931] = 36'h59350AF73;
        fsqrt_table[930] = 36'h590590F7B;
        fsqrt_table[929] = 36'h58D612F7E;
        fsqrt_table[928] = 36'h58A68AF87;
        fsqrt_table[927] = 36'h5876FEF8C;
        fsqrt_table[926] = 36'h58476AF93;
        fsqrt_table[925] = 36'h5817D0F9A;
        fsqrt_table[924] = 36'h57E830F9F;
        fsqrt_table[923] = 36'h57B888FA7;
        fsqrt_table[922] = 36'h5788DAFAD;
        fsqrt_table[921] = 36'h575926FB3;
        fsqrt_table[920] = 36'h57296AFBB;
        fsqrt_table[919] = 36'h56F9A8FC2;
        fsqrt_table[918] = 36'h56C9E0FC8;
        fsqrt_table[917] = 36'h569A10FD0;
        fsqrt_table[916] = 36'h566A3AFD7;
        fsqrt_table[915] = 36'h563A5EFDC;
        fsqrt_table[914] = 36'h560A7CFE1;
        fsqrt_table[913] = 36'h55DA92FE8;
        fsqrt_table[912] = 36'h55AAA0FF1;
        fsqrt_table[911] = 36'h557AA8FF9;
        fsqrt_table[910] = 36'h554AAAFFF;
        fsqrt_table[909] = 36'h551AA7004;
        fsqrt_table[908] = 36'h54EA9B00C;
        fsqrt_table[907] = 36'h54BA89012;
        fsqrt_table[906] = 36'h548A6F01A;
        fsqrt_table[905] = 36'h545A4F021;
        fsqrt_table[904] = 36'h542A29026;
        fsqrt_table[903] = 36'h53F9FB02E;
        fsqrt_table[902] = 36'h53C9C7034;
        fsqrt_table[901] = 36'h53998B03C;
        fsqrt_table[900] = 36'h536949042;
        fsqrt_table[899] = 36'h533901048;
        fsqrt_table[898] = 36'h5308B104F;
        fsqrt_table[897] = 36'h52D859058;
        fsqrt_table[896] = 36'h52A7FB05F;
        fsqrt_table[895] = 36'h527797065;
        fsqrt_table[894] = 36'h52472B06D;
        fsqrt_table[893] = 36'h5216B9073;
        fsqrt_table[892] = 36'h51E63F07B;
        fsqrt_table[891] = 36'h51B5BF081;
        fsqrt_table[890] = 36'h518539086;
        fsqrt_table[889] = 36'h5154A9090;
        fsqrt_table[888] = 36'h512415094;
        fsqrt_table[887] = 36'h50F37909B;
        fsqrt_table[886] = 36'h50C2D50A3;
        fsqrt_table[885] = 36'h50922B0AA;
        fsqrt_table[884] = 36'h5061790B2;
        fsqrt_table[883] = 36'h5030C10B8;
        fsqrt_table[882] = 36'h5000010C0;
        fsqrt_table[881] = 36'h4FCF3B0C6;
        fsqrt_table[880] = 36'h4F9E6D0CD;
        fsqrt_table[879] = 36'h4F6D990D3;
        fsqrt_table[878] = 36'h4F3CBD0DB;
        fsqrt_table[877] = 36'h4F0BD90E3;
        fsqrt_table[876] = 36'h4EDAEF0EA;
        fsqrt_table[875] = 36'h4EA9FF0F0;
        fsqrt_table[874] = 36'h4E79050F9;
        fsqrt_table[873] = 36'h4E4805101;
        fsqrt_table[872] = 36'h4E16FF107;
        fsqrt_table[871] = 36'h4DE5F110E;
        fsqrt_table[870] = 36'h4DB4DB116;
        fsqrt_table[869] = 36'h4D83BF11D;
        fsqrt_table[868] = 36'h4D529B125;
        fsqrt_table[867] = 36'h4D217112A;
        fsqrt_table[866] = 36'h4CF03F131;
        fsqrt_table[865] = 36'h4CBF05139;
        fsqrt_table[864] = 36'h4C8DC513F;
        fsqrt_table[863] = 36'h4C5C7D147;
        fsqrt_table[862] = 36'h4C2B2D14F;
        fsqrt_table[861] = 36'h4BF9D7155;
        fsqrt_table[860] = 36'h4BC87915C;
        fsqrt_table[859] = 36'h4B9713165;
        fsqrt_table[858] = 36'h4B65A516E;
        fsqrt_table[857] = 36'h4B3433172;
        fsqrt_table[856] = 36'h4B02B717A;
        fsqrt_table[855] = 36'h4AD133183;
        fsqrt_table[854] = 36'h4A9FA918A;
        fsqrt_table[853] = 36'h4A6E17192;
        fsqrt_table[852] = 36'h4A3C7F198;
        fsqrt_table[851] = 36'h4A0ADD1A1;
        fsqrt_table[850] = 36'h49D9351A9;
        fsqrt_table[849] = 36'h49A7851B1;
        fsqrt_table[848] = 36'h4975CF1B6;
        fsqrt_table[847] = 36'h4944111BD;
        fsqrt_table[846] = 36'h49124B1C4;
        fsqrt_table[845] = 36'h48E07D1CC;
        fsqrt_table[844] = 36'h48AEA71D5;
        fsqrt_table[843] = 36'h487CCB1DC;
        fsqrt_table[842] = 36'h484AE51E6;
        fsqrt_table[841] = 36'h4818FB1EA;
        fsqrt_table[840] = 36'h47E7071F3;
        fsqrt_table[839] = 36'h47B50B1FC;
        fsqrt_table[838] = 36'h478309202;
        fsqrt_table[837] = 36'h4750FF209;
        fsqrt_table[836] = 36'h471EED211;
        fsqrt_table[835] = 36'h46ECD3219;
        fsqrt_table[834] = 36'h46BAB1222;
        fsqrt_table[833] = 36'h468889228;
        fsqrt_table[832] = 36'h465657231;
        fsqrt_table[831] = 36'h46241F238;
        fsqrt_table[830] = 36'h45F1DF23F;
        fsqrt_table[829] = 36'h45BF97247;
        fsqrt_table[828] = 36'h458D4724F;
        fsqrt_table[827] = 36'h455AEF258;
        fsqrt_table[826] = 36'h45289125D;
        fsqrt_table[825] = 36'h44F629266;
        fsqrt_table[824] = 36'h44C3B9270;
        fsqrt_table[823] = 36'h449143276;
        fsqrt_table[822] = 36'h445EC527D;
        fsqrt_table[821] = 36'h442C3D287;
        fsqrt_table[820] = 36'h43F9AF28E;
        fsqrt_table[819] = 36'h43C719296;
        fsqrt_table[818] = 36'h43947B29D;
        fsqrt_table[817] = 36'h4361D52A5;
        fsqrt_table[816] = 36'h432F272AD;
        fsqrt_table[815] = 36'h42FC712B5;
        fsqrt_table[814] = 36'h42C9B32BD;
        fsqrt_table[813] = 36'h4296ED2C5;
        fsqrt_table[812] = 36'h42641F2CD;
        fsqrt_table[811] = 36'h4231492D5;
        fsqrt_table[810] = 36'h41FE6B2DD;
        fsqrt_table[809] = 36'h41CB852E5;
        fsqrt_table[808] = 36'h4198972ED;
        fsqrt_table[807] = 36'h4165A12F4;
        fsqrt_table[806] = 36'h4132A12FF;
        fsqrt_table[805] = 36'h40FF9B307;
        fsqrt_table[804] = 36'h40CC8D30E;
        fsqrt_table[803] = 36'h409977315;
        fsqrt_table[802] = 36'h40665731F;
        fsqrt_table[801] = 36'h403331326;
        fsqrt_table[800] = 36'h400001330;
        fsqrt_table[799] = 36'h3FCCCB336;
        fsqrt_table[798] = 36'h3F998B33F;
        fsqrt_table[797] = 36'h3F6643347;
        fsqrt_table[796] = 36'h3F32F3350;
        fsqrt_table[795] = 36'h3EFF9B358;
        fsqrt_table[794] = 36'h3ECC3B35F;
        fsqrt_table[793] = 36'h3E98D1369;
        fsqrt_table[792] = 36'h3E6561370;
        fsqrt_table[791] = 36'h3E31E7379;
        fsqrt_table[790] = 36'h3DFE65382;
        fsqrt_table[789] = 36'h3DCADB38A;
        fsqrt_table[788] = 36'h3D9749392;
        fsqrt_table[787] = 36'h3D63AF399;
        fsqrt_table[786] = 36'h3D300B3A3;
        fsqrt_table[785] = 36'h3CFC5F3AC;
        fsqrt_table[784] = 36'h3CC8AB3B4;
        fsqrt_table[783] = 36'h3C94EF3BC;
        fsqrt_table[782] = 36'h3C61293C6;
        fsqrt_table[781] = 36'h3C2D5D3CC;
        fsqrt_table[780] = 36'h3BF9873D5;
        fsqrt_table[779] = 36'h3BC5A93DC;
        fsqrt_table[778] = 36'h3B91C13E6;
        fsqrt_table[777] = 36'h3B5DD13F0;
        fsqrt_table[776] = 36'h3B29D93F8;
        fsqrt_table[775] = 36'h3AF5D9400;
        fsqrt_table[774] = 36'h3AC1CF40A;
        fsqrt_table[773] = 36'h3A8DBD413;
        fsqrt_table[772] = 36'h3A59A341A;
        fsqrt_table[771] = 36'h3A2581421;
        fsqrt_table[770] = 36'h39F15542A;
        fsqrt_table[769] = 36'h39BD21433;
        fsqrt_table[768] = 36'h3988E343C;
        fsqrt_table[767] = 36'h39549D445;
        fsqrt_table[766] = 36'h39204F44D;
        fsqrt_table[765] = 36'h38EBF7457;
        fsqrt_table[764] = 36'h38B797460;
        fsqrt_table[763] = 36'h38832F467;
        fsqrt_table[762] = 36'h384EBD471;
        fsqrt_table[761] = 36'h381A4147C;
        fsqrt_table[760] = 36'h37E5BF483;
        fsqrt_table[759] = 36'h37B13348B;
        fsqrt_table[758] = 36'h377C9D496;
        fsqrt_table[757] = 36'h3747FF49F;
        fsqrt_table[756] = 36'h3713594A7;
        fsqrt_table[755] = 36'h36DEA94B0;
        fsqrt_table[754] = 36'h36A9F14B8;
        fsqrt_table[753] = 36'h36752F4C1;
        fsqrt_table[752] = 36'h3640654CA;
        fsqrt_table[751] = 36'h360B914D3;
        fsqrt_table[750] = 36'h35D6B54DB;
        fsqrt_table[749] = 36'h35A1CF4E5;
        fsqrt_table[748] = 36'h356CE14ED;
        fsqrt_table[747] = 36'h3537E94F7;
        fsqrt_table[746] = 36'h3502E7502;
        fsqrt_table[745] = 36'h34CDDF508;
        fsqrt_table[744] = 36'h3498CB513;
        fsqrt_table[743] = 36'h3463AF51C;
        fsqrt_table[742] = 36'h342E89526;
        fsqrt_table[741] = 36'h33F95B52F;
        fsqrt_table[740] = 36'h33C425535;
        fsqrt_table[739] = 36'h338EE3540;
        fsqrt_table[738] = 36'h335999549;
        fsqrt_table[737] = 36'h332445554;
        fsqrt_table[736] = 36'h32EEE955C;
        fsqrt_table[735] = 36'h32B983566;
        fsqrt_table[734] = 36'h32841556D;
        fsqrt_table[733] = 36'h324E9B579;
        fsqrt_table[732] = 36'h32191B580;
        fsqrt_table[731] = 36'h31E38F58A;
        fsqrt_table[730] = 36'h31ADFB593;
        fsqrt_table[729] = 36'h31785D59C;
        fsqrt_table[728] = 36'h3142B55A6;
        fsqrt_table[727] = 36'h310D035B2;
        fsqrt_table[726] = 36'h30D7495BB;
        fsqrt_table[725] = 36'h30A1855C5;
        fsqrt_table[724] = 36'h306BB95CC;
        fsqrt_table[723] = 36'h3035E15D8;
        fsqrt_table[722] = 36'h3000015E1;
        fsqrt_table[721] = 36'h2FCA175EB;
        fsqrt_table[720] = 36'h2F94255F2;
        fsqrt_table[719] = 36'h2F5E275FD;
        fsqrt_table[718] = 36'h2F2821606;
        fsqrt_table[717] = 36'h2EF21160F;
        fsqrt_table[716] = 36'h2EBBF7619;
        fsqrt_table[715] = 36'h2E85D3623;
        fsqrt_table[714] = 36'h2E4FA562E;
        fsqrt_table[713] = 36'h2E196F636;
        fsqrt_table[712] = 36'h2DE32F63F;
        fsqrt_table[711] = 36'h2DACE364B;
        fsqrt_table[710] = 36'h2D7691652;
        fsqrt_table[709] = 36'h2D403165E;
        fsqrt_table[708] = 36'h2D09C9668;
        fsqrt_table[707] = 36'h2CD35966F;
        fsqrt_table[706] = 36'h2C9CDD67A;
        fsqrt_table[705] = 36'h2C6657685;
        fsqrt_table[704] = 36'h2C2FC968D;
        fsqrt_table[703] = 36'h2BF92F697;
        fsqrt_table[702] = 36'h2BC28B6A2;
        fsqrt_table[701] = 36'h2B8BDD6AE;
        fsqrt_table[700] = 36'h2B55276B6;
        fsqrt_table[699] = 36'h2B1E656C1;
        fsqrt_table[698] = 36'h2AE79B6C9;
        fsqrt_table[697] = 36'h2AB0C56D4;
        fsqrt_table[696] = 36'h2A79E56E0;
        fsqrt_table[695] = 36'h2A42FD6E7;
        fsqrt_table[694] = 36'h2A0C096F2;
        fsqrt_table[693] = 36'h29D50B6FD;
        fsqrt_table[692] = 36'h299E03707;
        fsqrt_table[691] = 36'h2966F1711;
        fsqrt_table[690] = 36'h292FD571B;
        fsqrt_table[689] = 36'h28F8AF725;
        fsqrt_table[688] = 36'h28C17D731;
        fsqrt_table[687] = 36'h288A4373A;
        fsqrt_table[686] = 36'h2852FD745;
        fsqrt_table[685] = 36'h281BAD750;
        fsqrt_table[684] = 36'h27E45375A;
        fsqrt_table[683] = 36'h27ACEF764;
        fsqrt_table[682] = 36'h27758176E;
        fsqrt_table[681] = 36'h273E07779;
        fsqrt_table[680] = 36'h270685781;
        fsqrt_table[679] = 36'h26CEF578F;
        fsqrt_table[678] = 36'h26975D799;
        fsqrt_table[677] = 36'h265FBB7A2;
        fsqrt_table[676] = 36'h26280D7AD;
        fsqrt_table[675] = 36'h25F0557B8;
        fsqrt_table[674] = 36'h25B8937C1;
        fsqrt_table[673] = 36'h2580C57CD;
        fsqrt_table[672] = 36'h2548ED7D8;
        fsqrt_table[671] = 36'h25110B7E2;
        fsqrt_table[670] = 36'h24D91D7EE;
        fsqrt_table[669] = 36'h24A1257F9;
        fsqrt_table[668] = 36'h246923803;
        fsqrt_table[667] = 36'h24311780C;
        fsqrt_table[666] = 36'h23F8FF816;
        fsqrt_table[665] = 36'h23C0DB823;
        fsqrt_table[664] = 36'h2388AF82B;
        fsqrt_table[663] = 36'h235075839;
        fsqrt_table[662] = 36'h231833842;
        fsqrt_table[661] = 36'h22DFE584C;
        fsqrt_table[660] = 36'h22A78B858;
        fsqrt_table[659] = 36'h226F27863;
        fsqrt_table[658] = 36'h2236B986D;
        fsqrt_table[657] = 36'h21FE3D87B;
        fsqrt_table[656] = 36'h21C5B9884;
        fsqrt_table[655] = 36'h218D2988F;
        fsqrt_table[654] = 36'h21548D89C;
        fsqrt_table[653] = 36'h211BE78A7;
        fsqrt_table[652] = 36'h20E3378B0;
        fsqrt_table[651] = 36'h20AA7B8BB;
        fsqrt_table[650] = 36'h2071B38C6;
        fsqrt_table[649] = 36'h2038E18D1;
        fsqrt_table[648] = 36'h2000018DF;
        fsqrt_table[647] = 36'h1FC7198E8;
        fsqrt_table[646] = 36'h1F8E258F3;
        fsqrt_table[645] = 36'h1F55258FF;
        fsqrt_table[644] = 36'h1F1C1B908;
        fsqrt_table[643] = 36'h1EE303916;
        fsqrt_table[642] = 36'h1EA9E1922;
        fsqrt_table[641] = 36'h1E70B592C;
        fsqrt_table[640] = 36'h1E377B939;
        fsqrt_table[639] = 36'h1DFE39942;
        fsqrt_table[638] = 36'h1DC4E994E;
        fsqrt_table[637] = 36'h1D8B8D95B;
        fsqrt_table[636] = 36'h1D5227965;
        fsqrt_table[635] = 36'h1D18B5971;
        fsqrt_table[634] = 36'h1CDF3797D;
        fsqrt_table[633] = 36'h1CA5AF987;
        fsqrt_table[632] = 36'h1C6C19994;
        fsqrt_table[631] = 36'h1C327999F;
        fsqrt_table[630] = 36'h1BF8CB9AD;
        fsqrt_table[629] = 36'h1BBF159B6;
        fsqrt_table[628] = 36'h1B85519C2;
        fsqrt_table[627] = 36'h1B4B819CE;
        fsqrt_table[626] = 36'h1B11A59DB;
        fsqrt_table[625] = 36'h1AD7BF9E5;
        fsqrt_table[624] = 36'h1A9DCB9F3;
        fsqrt_table[623] = 36'h1A63CD9FD;
        fsqrt_table[622] = 36'h1A29C1A0B;
        fsqrt_table[621] = 36'h19EFABA15;
        fsqrt_table[620] = 36'h19B587A23;
        fsqrt_table[619] = 36'h197B59A2E;
        fsqrt_table[618] = 36'h19411FA39;
        fsqrt_table[617] = 36'h1906D7A47;
        fsqrt_table[616] = 36'h18CC85A51;
        fsqrt_table[615] = 36'h189225A5F;
        fsqrt_table[614] = 36'h1857B9A6C;
        fsqrt_table[613] = 36'h181D43A76;
        fsqrt_table[612] = 36'h17E2BFA83;
        fsqrt_table[611] = 36'h17A82FA8F;
        fsqrt_table[610] = 36'h176D93A9B;
        fsqrt_table[609] = 36'h1732EBAA7;
        fsqrt_table[608] = 36'h16F835AB5;
        fsqrt_table[607] = 36'h16BD75ABF;
        fsqrt_table[606] = 36'h1682A7ACC;
        fsqrt_table[605] = 36'h1647CDAD9;
        fsqrt_table[604] = 36'h160CE7AE5;
        fsqrt_table[603] = 36'h15D1F3AF3;
        fsqrt_table[602] = 36'h1596F3B00;
        fsqrt_table[601] = 36'h155BE9B0A;
        fsqrt_table[600] = 36'h1520CFB18;
        fsqrt_table[599] = 36'h14E5ABB23;
        fsqrt_table[598] = 36'h14AA79B30;
        fsqrt_table[597] = 36'h146F39B3F;
        fsqrt_table[596] = 36'h1433EFB4A;
        fsqrt_table[595] = 36'h13F897B57;
        fsqrt_table[594] = 36'h13BD33B62;
        fsqrt_table[593] = 36'h1381C1B70;
        fsqrt_table[592] = 36'h134641B7F;
        fsqrt_table[591] = 36'h130AB7B8A;
        fsqrt_table[590] = 36'h12CF1FB97;
        fsqrt_table[589] = 36'h129379BA5;
        fsqrt_table[588] = 36'h1257C7BB2;
        fsqrt_table[587] = 36'h121C09BBD;
        fsqrt_table[586] = 36'h11E03DBCA;
        fsqrt_table[585] = 36'h11A463BD9;
        fsqrt_table[584] = 36'h11687DBE5;
        fsqrt_table[583] = 36'h112C89BF3;
        fsqrt_table[582] = 36'h10F089C00;
        fsqrt_table[581] = 36'h10B47BC0D;
        fsqrt_table[580] = 36'h107861C19;
        fsqrt_table[579] = 36'h103C39C26;
        fsqrt_table[578] = 36'h100003C34;
        fsqrt_table[577] = 36'h0FC3BFC43;
        fsqrt_table[576] = 36'h0F876FC50;
        fsqrt_table[575] = 36'h0F4B13C5B;
        fsqrt_table[574] = 36'h0F0EA7C69;
        fsqrt_table[573] = 36'h0ED22DC79;
        fsqrt_table[572] = 36'h0E95A7C86;
        fsqrt_table[571] = 36'h0E5915C91;
        fsqrt_table[570] = 36'h0E1C73CA0;
        fsqrt_table[569] = 36'h0DDFC5CAC;
        fsqrt_table[568] = 36'h0DA307CBC;
        fsqrt_table[567] = 36'h0D663DCC9;
        fsqrt_table[566] = 36'h0D2965CD7;
        fsqrt_table[565] = 36'h0CEC7FCE6;
        fsqrt_table[564] = 36'h0CAF8BCF4;
        fsqrt_table[563] = 36'h0C728BD00;
        fsqrt_table[562] = 36'h0C357BD0F;
        fsqrt_table[561] = 36'h0BF85FD1B;
        fsqrt_table[560] = 36'h0BBB33D2A;
        fsqrt_table[559] = 36'h0B7DFBD37;
        fsqrt_table[558] = 36'h0B40B3D46;
        fsqrt_table[557] = 36'h0B035DD55;
        fsqrt_table[556] = 36'h0AC5FBD61;
        fsqrt_table[555] = 36'h0A8889D70;
        fsqrt_table[554] = 36'h0A4B09D7F;
        fsqrt_table[553] = 36'h0A0D7BD8E;
        fsqrt_table[552] = 36'h09CFDFD9C;
        fsqrt_table[551] = 36'h099235DAA;
        fsqrt_table[550] = 36'h09547DDB7;
        fsqrt_table[549] = 36'h0916B5DC7;
        fsqrt_table[548] = 36'h08D8E1DD3;
        fsqrt_table[547] = 36'h089AFDDE1;
        fsqrt_table[546] = 36'h085D09DF2;
        fsqrt_table[545] = 36'h081F09DFF;
        fsqrt_table[544] = 36'h07E0F9E0F;
        fsqrt_table[543] = 36'h07A2DBE1D;
        fsqrt_table[542] = 36'h0764AFE2A;
        fsqrt_table[541] = 36'h072673E3A;
        fsqrt_table[540] = 36'h06E829E48;
        fsqrt_table[539] = 36'h06A9CFE59;
        fsqrt_table[538] = 36'h066B69E65;
        fsqrt_table[537] = 36'h062CF1E76;
        fsqrt_table[536] = 36'h05EE6BE86;
        fsqrt_table[535] = 36'h05AFD7E94;
        fsqrt_table[534] = 36'h057135EA1;
        fsqrt_table[533] = 36'h053281EB2;
        fsqrt_table[532] = 36'h04F3C1EBF;
        fsqrt_table[531] = 36'h04B4EFED0;
        fsqrt_table[530] = 36'h04760FEDF;
        fsqrt_table[529] = 36'h043721EED;
        fsqrt_table[528] = 36'h03F823EFC;
        fsqrt_table[527] = 36'h03B915F0C;
        fsqrt_table[526] = 36'h0379F9F1A;
        fsqrt_table[525] = 36'h033ACBF2C;
        fsqrt_table[524] = 36'h02FB91F39;
        fsqrt_table[523] = 36'h02BC45F4A;
        fsqrt_table[522] = 36'h027CEBF59;
        fsqrt_table[521] = 36'h023D81F68;
        fsqrt_table[520] = 36'h01FE07F78;
        fsqrt_table[519] = 36'h01BE7DF89;
        fsqrt_table[518] = 36'h017EE5F97;
        fsqrt_table[517] = 36'h013F3BFA9;
        fsqrt_table[516] = 36'h00FF83FB8;
        fsqrt_table[515] = 36'h00BFBBFC7;
        fsqrt_table[514] = 36'h007FE3FD7;
        fsqrt_table[513] = 36'h003FFBFE7;
        fsqrt_table[512] = 36'h000003FF7;
        fsqrt_table[511] = 36'hFFBFFC002;
        fsqrt_table[510] = 36'hFF7FF0006;
        fsqrt_table[509] = 36'hFF3FDC00A;
        fsqrt_table[508] = 36'hFEFFC000E;
        fsqrt_table[507] = 36'hFEBF9C012;
        fsqrt_table[506] = 36'hFE7F70016;
        fsqrt_table[505] = 36'hFE3F3C01A;
        fsqrt_table[504] = 36'hFDFF0001E;
        fsqrt_table[503] = 36'hFDBEBA023;
        fsqrt_table[502] = 36'hFD7E70025;
        fsqrt_table[501] = 36'hFD3E1A02A;
        fsqrt_table[500] = 36'hFCFDBE02E;
        fsqrt_table[499] = 36'hFCBD5A031;
        fsqrt_table[498] = 36'hFC7CEC036;
        fsqrt_table[497] = 36'hFC3C78039;
        fsqrt_table[496] = 36'hFBFBF803F;
        fsqrt_table[495] = 36'hFBBB74042;
        fsqrt_table[494] = 36'hFB7AE6046;
        fsqrt_table[493] = 36'hFB3A5004A;
        fsqrt_table[492] = 36'hFAF9B204E;
        fsqrt_table[491] = 36'hFAB90A053;
        fsqrt_table[490] = 36'hFA785C057;
        fsqrt_table[489] = 36'hFA37A605A;
        fsqrt_table[488] = 36'hF9F6E605F;
        fsqrt_table[487] = 36'hF9B61E063;
        fsqrt_table[486] = 36'hF9754E068;
        fsqrt_table[485] = 36'hF9347606C;
        fsqrt_table[484] = 36'hF8F396070;
        fsqrt_table[483] = 36'hF8B2AE073;
        fsqrt_table[482] = 36'hF871BA079;
        fsqrt_table[481] = 36'hF830C207C;
        fsqrt_table[480] = 36'hF7EFC0080;
        fsqrt_table[479] = 36'hF7AEB6084;
        fsqrt_table[478] = 36'hF76DA4088;
        fsqrt_table[477] = 36'hF72C8808D;
        fsqrt_table[476] = 36'hF6EB64091;
        fsqrt_table[475] = 36'hF6AA38096;
        fsqrt_table[474] = 36'hF66904099;
        fsqrt_table[473] = 36'hF627C609E;
        fsqrt_table[472] = 36'hF5E6800A3;
        fsqrt_table[471] = 36'hF5A5320A7;
        fsqrt_table[470] = 36'hF563DC0AB;
        fsqrt_table[469] = 36'hF5227E0AF;
        fsqrt_table[468] = 36'hF4E1160B3;
        fsqrt_table[467] = 36'hF49FA60B8;
        fsqrt_table[466] = 36'hF45E2C0BD;
        fsqrt_table[465] = 36'hF41CAC0C0;
        fsqrt_table[464] = 36'hF3DB220C5;
        fsqrt_table[463] = 36'hF399900C9;
        fsqrt_table[462] = 36'hF357F40CE;
        fsqrt_table[461] = 36'hF316520D1;
        fsqrt_table[460] = 36'hF2D4A60D5;
        fsqrt_table[459] = 36'hF292F20D9;
        fsqrt_table[458] = 36'hF251320DF;
        fsqrt_table[457] = 36'hF20F6C0E3;
        fsqrt_table[456] = 36'hF1CD9E0E7;
        fsqrt_table[455] = 36'hF18BC80EA;
        fsqrt_table[454] = 36'hF149E60F0;
        fsqrt_table[453] = 36'hF107FE0F3;
        fsqrt_table[452] = 36'hF0C60C0F8;
        fsqrt_table[451] = 36'hF084100FD;
        fsqrt_table[450] = 36'hF0420C102;
        fsqrt_table[449] = 36'hF00002105;
        fsqrt_table[448] = 36'hEFBDEC10A;
        fsqrt_table[447] = 36'hEF7BCE10F;
        fsqrt_table[446] = 36'hEF39A8113;
        fsqrt_table[445] = 36'hEEF77A116;
        fsqrt_table[444] = 36'hEEB54011C;
        fsqrt_table[443] = 36'hEE72FE121;
        fsqrt_table[442] = 36'hEE30B6124;
        fsqrt_table[441] = 36'hEDEE62129;
        fsqrt_table[440] = 36'hEDAC0612E;
        fsqrt_table[439] = 36'hED69A2132;
        fsqrt_table[438] = 36'hED2734136;
        fsqrt_table[437] = 36'hECE4BE13B;
        fsqrt_table[436] = 36'hECA23E13F;
        fsqrt_table[435] = 36'hEC5FB6143;
        fsqrt_table[434] = 36'hEC1D24148;
        fsqrt_table[433] = 36'hEBDA8A14C;
        fsqrt_table[432] = 36'hEB97E6151;
        fsqrt_table[431] = 36'hEB553A155;
        fsqrt_table[430] = 36'hEB128215B;
        fsqrt_table[429] = 36'hEACFC415F;
        fsqrt_table[428] = 36'hEA8CFC164;
        fsqrt_table[427] = 36'hEA4A2C168;
        fsqrt_table[426] = 36'hEA075216C;
        fsqrt_table[425] = 36'hE9C470170;
        fsqrt_table[424] = 36'hE98182176;
        fsqrt_table[423] = 36'hE93E8E179;
        fsqrt_table[422] = 36'hE8FB8E17F;
        fsqrt_table[421] = 36'hE8B886184;
        fsqrt_table[420] = 36'hE87574189;
        fsqrt_table[419] = 36'hE8325A18D;
        fsqrt_table[418] = 36'hE7EF38191;
        fsqrt_table[417] = 36'hE7AC0C195;
        fsqrt_table[416] = 36'hE768D419B;
        fsqrt_table[415] = 36'hE7259619F;
        fsqrt_table[414] = 36'hE6E24E1A3;
        fsqrt_table[413] = 36'hE69EFC1A8;
        fsqrt_table[412] = 36'hE65BA01AD;
        fsqrt_table[411] = 36'hE6183C1B2;
        fsqrt_table[410] = 36'hE5D4CE1B6;
        fsqrt_table[409] = 36'hE591581BA;
        fsqrt_table[408] = 36'hE54DD61C0;
        fsqrt_table[407] = 36'hE50A4C1C5;
        fsqrt_table[406] = 36'hE4C6BA1C8;
        fsqrt_table[405] = 36'hE4831C1CE;
        fsqrt_table[404] = 36'hE43F761D2;
        fsqrt_table[403] = 36'hE3FBC61D7;
        fsqrt_table[402] = 36'hE3B80E1DB;
        fsqrt_table[401] = 36'hE3744A1E1;
        fsqrt_table[400] = 36'hE3307E1E6;
        fsqrt_table[399] = 36'hE2ECAA1E9;
        fsqrt_table[398] = 36'hE2A8C81F0;
        fsqrt_table[397] = 36'hE264E01F4;
        fsqrt_table[396] = 36'hE220EE1F9;
        fsqrt_table[395] = 36'hE1DCF21FE;
        fsqrt_table[394] = 36'hE198EE202;
        fsqrt_table[393] = 36'hE154DE207;
        fsqrt_table[392] = 36'hE110C620B;
        fsqrt_table[391] = 36'hE0CCA2211;
        fsqrt_table[390] = 36'hE08876216;
        fsqrt_table[389] = 36'hE0444021B;
        fsqrt_table[388] = 36'hE00000220;
        fsqrt_table[387] = 36'hDFBBB8224;
        fsqrt_table[386] = 36'hDF7766229;
        fsqrt_table[385] = 36'hDF330822E;
        fsqrt_table[384] = 36'hDEEEA2233;
        fsqrt_table[383] = 36'hDEAA32238;
        fsqrt_table[382] = 36'hDE65B823D;
        fsqrt_table[381] = 36'hDE2134242;
        fsqrt_table[380] = 36'hDDDCA6247;
        fsqrt_table[379] = 36'hDD981024B;
        fsqrt_table[378] = 36'hDD537024F;
        fsqrt_table[377] = 36'hDD0EC2256;
        fsqrt_table[376] = 36'hDCCA0E25A;
        fsqrt_table[375] = 36'hDC854E260;
        fsqrt_table[374] = 36'hDC4086264;
        fsqrt_table[373] = 36'hDBFBB4269;
        fsqrt_table[372] = 36'hDBB6D826D;
        fsqrt_table[371] = 36'hDB71F0273;
        fsqrt_table[370] = 36'hDB2D00278;
        fsqrt_table[369] = 36'hDAE80627C;
        fsqrt_table[368] = 36'hDAA300282;
        fsqrt_table[367] = 36'hDA5DF0288;
        fsqrt_table[366] = 36'hDA18DA28B;
        fsqrt_table[365] = 36'hD9D3B6291;
        fsqrt_table[364] = 36'hD98E8A295;
        fsqrt_table[363] = 36'hD9495229B;
        fsqrt_table[362] = 36'hD9041229F;
        fsqrt_table[361] = 36'hD8BEC42A6;
        fsqrt_table[360] = 36'hD879702AA;
        fsqrt_table[359] = 36'hD834102AF;
        fsqrt_table[358] = 36'hD7EEA62B4;
        fsqrt_table[357] = 36'hD7A9322B9;
        fsqrt_table[356] = 36'hD763B42BE;
        fsqrt_table[355] = 36'hD71E2C2C3;
        fsqrt_table[354] = 36'hD6D8982C9;
        fsqrt_table[353] = 36'hD692FC2CD;
        fsqrt_table[352] = 36'hD64D522D4;
        fsqrt_table[351] = 36'hD607A22D8;
        fsqrt_table[350] = 36'hD5C1E62DD;
        fsqrt_table[349] = 36'hD57C1E2E3;
        fsqrt_table[348] = 36'hD5364E2E8;
        fsqrt_table[347] = 36'hD4F0742EC;
        fsqrt_table[346] = 36'hD4AA8C2F3;
        fsqrt_table[345] = 36'hD4649C2F8;
        fsqrt_table[344] = 36'hD41EA22FD;
        fsqrt_table[343] = 36'hD3D89E302;
        fsqrt_table[342] = 36'hD3928E307;
        fsqrt_table[341] = 36'hD34C7430C;
        fsqrt_table[340] = 36'hD30650311;
        fsqrt_table[339] = 36'hD2C020317;
        fsqrt_table[338] = 36'hD279E831B;
        fsqrt_table[337] = 36'hD233A2322;
        fsqrt_table[336] = 36'hD1ED54327;
        fsqrt_table[335] = 36'hD1A6FA32C;
        fsqrt_table[334] = 36'hD16096332;
        fsqrt_table[333] = 36'hD11A28336;
        fsqrt_table[332] = 36'hD0D3AE33C;
        fsqrt_table[331] = 36'hD08D2A341;
        fsqrt_table[330] = 36'hD0469C346;
        fsqrt_table[329] = 36'hD0000234C;
        fsqrt_table[328] = 36'hCFB95E351;
        fsqrt_table[327] = 36'hCF72AE357;
        fsqrt_table[326] = 36'hCF2BF435D;
        fsqrt_table[325] = 36'hCEE530362;
        fsqrt_table[324] = 36'hCE9E60367;
        fsqrt_table[323] = 36'hCE578636D;
        fsqrt_table[322] = 36'hCE10A2371;
        fsqrt_table[321] = 36'hCDC9B0378;
        fsqrt_table[320] = 36'hCD82B637D;
        fsqrt_table[319] = 36'hCD3BB0382;
        fsqrt_table[318] = 36'hCCF4A0387;
        fsqrt_table[317] = 36'hCCAD8438D;
        fsqrt_table[316] = 36'hCC665C393;
        fsqrt_table[315] = 36'hCC1F2A399;
        fsqrt_table[314] = 36'hCBD7EE39E;
        fsqrt_table[313] = 36'hCB90A63A4;
        fsqrt_table[312] = 36'hCB49543A8;
        fsqrt_table[311] = 36'hCB01F63AE;
        fsqrt_table[310] = 36'hCABA8C3B4;
        fsqrt_table[309] = 36'hCA73183BA;
        fsqrt_table[308] = 36'hCA2B9A3BE;
        fsqrt_table[307] = 36'hC9E40E3C5;
        fsqrt_table[306] = 36'hC99C783CB;
        fsqrt_table[305] = 36'hC954D83D0;
        fsqrt_table[304] = 36'hC90D2C3D5;
        fsqrt_table[303] = 36'hC8C5743DB;
        fsqrt_table[302] = 36'hC87DB23E0;
        fsqrt_table[301] = 36'hC835E43E6;
        fsqrt_table[300] = 36'hC7EE0A3EC;
        fsqrt_table[299] = 36'hC7A6263F2;
        fsqrt_table[298] = 36'hC75E363F7;
        fsqrt_table[297] = 36'hC7163A3FD;
        fsqrt_table[296] = 36'hC6CE34403;
        fsqrt_table[295] = 36'hC68622408;
        fsqrt_table[294] = 36'hC63E0440E;
        fsqrt_table[293] = 36'hC5F5DC413;
        fsqrt_table[292] = 36'hC5ADA641A;
        fsqrt_table[291] = 36'hC56566420;
        fsqrt_table[290] = 36'hC51D1A426;
        fsqrt_table[289] = 36'hC4D4C442B;
        fsqrt_table[288] = 36'hC48C62431;
        fsqrt_table[287] = 36'hC443F4436;
        fsqrt_table[286] = 36'hC3FB7A43C;
        fsqrt_table[285] = 36'hC3B2F4442;
        fsqrt_table[284] = 36'hC36A64447;
        fsqrt_table[283] = 36'hC321C644E;
        fsqrt_table[282] = 36'hC2D91E454;
        fsqrt_table[281] = 36'hC2906A459;
        fsqrt_table[280] = 36'hC247AA45F;
        fsqrt_table[279] = 36'hC1FEDE466;
        fsqrt_table[278] = 36'hC1B60846A;
        fsqrt_table[277] = 36'hC16D24471;
        fsqrt_table[276] = 36'hC12434478;
        fsqrt_table[275] = 36'hC0DB3A47D;
        fsqrt_table[274] = 36'hC09234482;
        fsqrt_table[273] = 36'hC04920489;
        fsqrt_table[272] = 36'hC0000248F;
        fsqrt_table[271] = 36'hBFB6D8494;
        fsqrt_table[270] = 36'hBF6DA049B;
        fsqrt_table[269] = 36'hBF245E4A1;
        fsqrt_table[268] = 36'hBEDB104A6;
        fsqrt_table[267] = 36'hBE91B64AC;
        fsqrt_table[266] = 36'hBE484E4B3;
        fsqrt_table[265] = 36'hBDFEDC4B9;
        fsqrt_table[264] = 36'hBDB55E4BE;
        fsqrt_table[263] = 36'hBD6BD24C5;
        fsqrt_table[262] = 36'hBD223C4CA;
        fsqrt_table[261] = 36'hBCD8984D1;
        fsqrt_table[260] = 36'hBC8EE84D8;
        fsqrt_table[259] = 36'hBC452E4DC;
        fsqrt_table[258] = 36'hBBFB644E4;
        fsqrt_table[257] = 36'hBBB1904EA;
        fsqrt_table[256] = 36'hBB67B04F0;
        fsqrt_table[255] = 36'hBB1DC44F5;
        fsqrt_table[254] = 36'hBAD3CA4FC;
        fsqrt_table[253] = 36'hBA89C6501;
        fsqrt_table[252] = 36'hBA3FB2509;
        fsqrt_table[251] = 36'hB9F59450F;
        fsqrt_table[250] = 36'hB9AB6A515;
        fsqrt_table[249] = 36'hB9613451A;
        fsqrt_table[248] = 36'hB916EE522;
        fsqrt_table[247] = 36'hB8CC9E528;
        fsqrt_table[246] = 36'hB8824252E;
        fsqrt_table[245] = 36'hB837DA533;
        fsqrt_table[244] = 36'hB7ED6253B;
        fsqrt_table[243] = 36'hB7A2E0541;
        fsqrt_table[242] = 36'hB75852547;
        fsqrt_table[241] = 36'hB70DB654D;
        fsqrt_table[240] = 36'hB6C30E553;
        fsqrt_table[239] = 36'hB6785855A;
        fsqrt_table[238] = 36'hB62D96561;
        fsqrt_table[237] = 36'hB5E2C8566;
        fsqrt_table[236] = 36'hB597EC56D;
        fsqrt_table[235] = 36'hB54D04573;
        fsqrt_table[234] = 36'hB5020E57B;
        fsqrt_table[233] = 36'hB4B70C581;
        fsqrt_table[232] = 36'hB46BFE587;
        fsqrt_table[231] = 36'hB420E258D;
        fsqrt_table[230] = 36'hB3D5BA593;
        fsqrt_table[229] = 36'hB38A8459A;
        fsqrt_table[228] = 36'hB33F425A0;
        fsqrt_table[227] = 36'hB2F3F05A8;
        fsqrt_table[226] = 36'hB2A8945AE;
        fsqrt_table[225] = 36'hB25D2A5B5;
        fsqrt_table[224] = 36'hB211B45BB;
        fsqrt_table[223] = 36'hB1C6305C1;
        fsqrt_table[222] = 36'hB17A9E5C8;
        fsqrt_table[221] = 36'hB12F005CF;
        fsqrt_table[220] = 36'hB0E3545D5;
        fsqrt_table[219] = 36'hB0979C5DB;
        fsqrt_table[218] = 36'hB04BD65E2;
        fsqrt_table[217] = 36'hB000025E9;
        fsqrt_table[216] = 36'hAFB4225EF;
        fsqrt_table[215] = 36'hAF68325F7;
        fsqrt_table[214] = 36'hAF1C385FD;
        fsqrt_table[213] = 36'hAED02E604;
        fsqrt_table[212] = 36'hAE841860B;
        fsqrt_table[211] = 36'hAE37F4612;
        fsqrt_table[210] = 36'hADEBC4618;
        fsqrt_table[209] = 36'hAD9F8461F;
        fsqrt_table[208] = 36'hAD5338626;
        fsqrt_table[207] = 36'hAD06DE62D;
        fsqrt_table[206] = 36'hACBA78633;
        fsqrt_table[205] = 36'hAC6E0263A;
        fsqrt_table[204] = 36'hAC2180640;
        fsqrt_table[203] = 36'hABD4F0647;
        fsqrt_table[202] = 36'hAB885064F;
        fsqrt_table[201] = 36'hAB3BA6655;
        fsqrt_table[200] = 36'hAAEEEC65C;
        fsqrt_table[199] = 36'hAAA224663;
        fsqrt_table[198] = 36'hAA554E66B;
        fsqrt_table[197] = 36'hAA086C671;
        fsqrt_table[196] = 36'hA9BB7A678;
        fsqrt_table[195] = 36'hA96E7C67F;
        fsqrt_table[194] = 36'hA9216E687;
        fsqrt_table[193] = 36'hA8D45468D;
        fsqrt_table[192] = 36'hA8872C693;
        fsqrt_table[191] = 36'hA839F469B;
        fsqrt_table[190] = 36'hA7ECB06A1;
        fsqrt_table[189] = 36'hA79F5C6A9;
        fsqrt_table[188] = 36'hA751FC6AF;
        fsqrt_table[187] = 36'hA7048C6B7;
        fsqrt_table[186] = 36'hA6B70E6BF;
        fsqrt_table[185] = 36'hA669826C6;
        fsqrt_table[184] = 36'hA61BE86CD;
        fsqrt_table[183] = 36'hA5CE406D4;
        fsqrt_table[182] = 36'hA5808A6DB;
        fsqrt_table[181] = 36'hA532C66E1;
        fsqrt_table[180] = 36'hA4E4F26E9;
        fsqrt_table[179] = 36'hA497106F0;
        fsqrt_table[178] = 36'hA449206F8;
        fsqrt_table[177] = 36'hA3FB226FE;
        fsqrt_table[176] = 36'hA3AD14706;
        fsqrt_table[175] = 36'hA35EFA70D;
        fsqrt_table[174] = 36'hA310CE715;
        fsqrt_table[173] = 36'hA2C29671C;
        fsqrt_table[172] = 36'hA2744E724;
        fsqrt_table[171] = 36'hA225F872B;
        fsqrt_table[170] = 36'hA1D794732;
        fsqrt_table[169] = 36'hA1892073A;
        fsqrt_table[168] = 36'hA13A9E741;
        fsqrt_table[167] = 36'hA0EC0E748;
        fsqrt_table[166] = 36'hA09D6E74F;
        fsqrt_table[165] = 36'hA04EC0756;
        fsqrt_table[164] = 36'hA0000275E;
        fsqrt_table[163] = 36'h9FB136765;
        fsqrt_table[162] = 36'h9F625A76D;
        fsqrt_table[161] = 36'h9F1370775;
        fsqrt_table[160] = 36'h9EC47677D;
        fsqrt_table[159] = 36'h9E756E784;
        fsqrt_table[158] = 36'h9E265678C;
        fsqrt_table[157] = 36'h9DD730793;
        fsqrt_table[156] = 36'h9D87FA79B;
        fsqrt_table[155] = 36'h9D38B67A2;
        fsqrt_table[154] = 36'h9CE9627A9;
        fsqrt_table[153] = 36'h9C99FE7B1;
        fsqrt_table[152] = 36'h9C4A8C7B8;
        fsqrt_table[151] = 36'h9BFB0A7C0;
        fsqrt_table[150] = 36'h9BAB787C8;
        fsqrt_table[149] = 36'h9B5BD87CF;
        fsqrt_table[148] = 36'h9B0C287D7;
        fsqrt_table[147] = 36'h9ABC687DF;
        fsqrt_table[146] = 36'h9A6C987E7;
        fsqrt_table[145] = 36'h9A1CBA7EF;
        fsqrt_table[144] = 36'h99CCCC7F6;
        fsqrt_table[143] = 36'h997CCE7FE;
        fsqrt_table[142] = 36'h992CC0807;
        fsqrt_table[141] = 36'h98DCA480E;
        fsqrt_table[140] = 36'h988C76816;
        fsqrt_table[139] = 36'h983C3A81E;
        fsqrt_table[138] = 36'h97EBEE825;
        fsqrt_table[137] = 36'h979B9282D;
        fsqrt_table[136] = 36'h974B26835;
        fsqrt_table[135] = 36'h96FAAA83D;
        fsqrt_table[134] = 36'h96AA1E845;
        fsqrt_table[133] = 36'h96598284D;
        fsqrt_table[132] = 36'h9608D6855;
        fsqrt_table[131] = 36'h95B81A85D;
        fsqrt_table[130] = 36'h95674E866;
        fsqrt_table[129] = 36'h95167286E;
        fsqrt_table[128] = 36'h94C586875;
        fsqrt_table[127] = 36'h94748A87D;
        fsqrt_table[126] = 36'h94237C886;
        fsqrt_table[125] = 36'h93D26088E;
        fsqrt_table[124] = 36'h938132897;
        fsqrt_table[123] = 36'h932FF489F;
        fsqrt_table[122] = 36'h92DEA88A6;
        fsqrt_table[121] = 36'h928D488AF;
        fsqrt_table[120] = 36'h923BDA8B7;
        fsqrt_table[119] = 36'h91EA5A8C0;
        fsqrt_table[118] = 36'h9198CA8C8;
        fsqrt_table[117] = 36'h91472A8D0;
        fsqrt_table[116] = 36'h90F57A8D8;
        fsqrt_table[115] = 36'h90A3B88E0;
        fsqrt_table[114] = 36'h9051E68E8;
        fsqrt_table[113] = 36'h9000028F1;
        fsqrt_table[112] = 36'h8FAE0E8FA;
        fsqrt_table[111] = 36'h8F5C0A902;
        fsqrt_table[110] = 36'h8F09F490A;
        fsqrt_table[109] = 36'h8EB7CE912;
        fsqrt_table[108] = 36'h8E659691B;
        fsqrt_table[107] = 36'h8E134E923;
        fsqrt_table[106] = 36'h8DC0F492C;
        fsqrt_table[105] = 36'h8D6E8A935;
        fsqrt_table[104] = 36'h8D1C0E93D;
        fsqrt_table[103] = 36'h8CC982945;
        fsqrt_table[102] = 36'h8C76E494E;
        fsqrt_table[101] = 36'h8C2434957;
        fsqrt_table[100] = 36'h8BD174960;
        fsqrt_table[99] = 36'h8B7EA2969;
        fsqrt_table[98] = 36'h8B2BBE972;
        fsqrt_table[97] = 36'h8AD8CA97A;
        fsqrt_table[96] = 36'h8A85C4983;
        fsqrt_table[95] = 36'h8A32AC98C;
        fsqrt_table[94] = 36'h89DF84994;
        fsqrt_table[93] = 36'h898C4A99D;
        fsqrt_table[92] = 36'h8938FE9A5;
        fsqrt_table[91] = 36'h88E5A09AE;
        fsqrt_table[90] = 36'h8892309B7;
        fsqrt_table[89] = 36'h883EAE9C1;
        fsqrt_table[88] = 36'h87EB1C9C9;
        fsqrt_table[87] = 36'h8797769D3;
        fsqrt_table[86] = 36'h8743C09DB;
        fsqrt_table[85] = 36'h86EFF89E3;
        fsqrt_table[84] = 36'h869C1C9EE;
        fsqrt_table[83] = 36'h8648309F6;
        fsqrt_table[82] = 36'h85F4329FE;
        fsqrt_table[81] = 36'h85A020A08;
        fsqrt_table[80] = 36'h854BFEA11;
        fsqrt_table[79] = 36'h84F7C8A1A;
        fsqrt_table[78] = 36'h84A380A24;
        fsqrt_table[77] = 36'h844F26A2D;
        fsqrt_table[76] = 36'h83FABAA35;
        fsqrt_table[75] = 36'h83A63CA3F;
        fsqrt_table[74] = 36'h8351ACA48;
        fsqrt_table[73] = 36'h82FD08A51;
        fsqrt_table[72] = 36'h82A852A5B;
        fsqrt_table[71] = 36'h82538AA64;
        fsqrt_table[70] = 36'h81FEAEA6E;
        fsqrt_table[69] = 36'h81A9C0A77;
        fsqrt_table[68] = 36'h8154C0A80;
        fsqrt_table[67] = 36'h80FFACA8A;
        fsqrt_table[66] = 36'h80AA86A92;
        fsqrt_table[65] = 36'h80554EA9C;
        fsqrt_table[64] = 36'h800002AA6;
        fsqrt_table[63] = 36'h7FAAA4AAF;
        fsqrt_table[62] = 36'h7F5532AB8;
        fsqrt_table[61] = 36'h7EFFACAC3;
        fsqrt_table[60] = 36'h7EAA14ACC;
        fsqrt_table[59] = 36'h7E546AAD5;
        fsqrt_table[58] = 36'h7DFEAAAE0;
        fsqrt_table[57] = 36'h7DA8DAAE8;
        fsqrt_table[56] = 36'h7D52F4AF3;
        fsqrt_table[55] = 36'h7CFCFCAFC;
        fsqrt_table[54] = 36'h7CA6F0B06;
        fsqrt_table[53] = 36'h7C50D0B0F;
        fsqrt_table[52] = 36'h7BFA9EB1A;
        fsqrt_table[51] = 36'h7BA458B23;
        fsqrt_table[50] = 36'h7B4DFEB2D;
        fsqrt_table[49] = 36'h7AF790B37;
        fsqrt_table[48] = 36'h7AA110B40;
        fsqrt_table[47] = 36'h7A4A7AB4B;
        fsqrt_table[46] = 36'h79F3D2B54;
        fsqrt_table[45] = 36'h799D14B5F;
        fsqrt_table[44] = 36'h794644B68;
        fsqrt_table[43] = 36'h78EF5EB73;
        fsqrt_table[42] = 36'h789866B7C;
        fsqrt_table[41] = 36'h784158B87;
        fsqrt_table[40] = 36'h77EA38B90;
        fsqrt_table[39] = 36'h779302B9B;
        fsqrt_table[38] = 36'h773BB8BA4;
        fsqrt_table[37] = 36'h76E45CBAE;
        fsqrt_table[36] = 36'h768CE8BBA;
        fsqrt_table[35] = 36'h763562BC2;
        fsqrt_table[34] = 36'h75DDC6BCD;
        fsqrt_table[33] = 36'h758618BD7;
        fsqrt_table[32] = 36'h752E52BE3;
        fsqrt_table[31] = 36'h74D67ABEC;
        fsqrt_table[30] = 36'h747E8CBF7;
        fsqrt_table[29] = 36'h74268AC01;
        fsqrt_table[28] = 36'h73CE72C0C;
        fsqrt_table[27] = 36'h737646C16;
        fsqrt_table[26] = 36'h731E04C20;
        fsqrt_table[25] = 36'h72C5AEC2A;
        fsqrt_table[24] = 36'h726D44C35;
        fsqrt_table[23] = 36'h7214C4C40;
        fsqrt_table[22] = 36'h71BC2EC4B;
        fsqrt_table[21] = 36'h716382C56;
        fsqrt_table[20] = 36'h710AC2C5F;
        fsqrt_table[19] = 36'h70B1EEC6A;
        fsqrt_table[18] = 36'h705902C76;
        fsqrt_table[17] = 36'h700002C80;
        fsqrt_table[16] = 36'h6FA6ECC8B;
        fsqrt_table[15] = 36'h6F4DC0C95;
        fsqrt_table[14] = 36'h6EF480CA0;
        fsqrt_table[13] = 36'h6E9B28CAC;
        fsqrt_table[12] = 36'h6E41BCCB6;
        fsqrt_table[11] = 36'h6DE83ACC1;
        fsqrt_table[10] = 36'h6D8EA0CCD;
        fsqrt_table[9] = 36'h6D34F2CD6;
        fsqrt_table[8] = 36'h6CDB2ECE2;
        fsqrt_table[7] = 36'h6C8154CED;
        fsqrt_table[6] = 36'h6C2762CF9;
        fsqrt_table[5] = 36'h6BCD5CD03;
        fsqrt_table[4] = 36'h6B733ED0F;
        fsqrt_table[3] = 36'h6B190AD1A;
        fsqrt_table[2] = 36'h6ABEC0D24;
        fsqrt_table[1] = 36'h6A6460D30;
        fsqrt_table[0] = 36'h6A09E8D3C;
    end

    always @(posedge clk) begin
        if (en) begin
            if (we)
                fsqrt_table[addr] <= di;
            if (rst)
                dout <= 0;
            else
                dout <= fsqrt_table[addr];
        end
    end

endmodule

`default_nettype wire