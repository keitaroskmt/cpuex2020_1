`default_nettype none

module finv
    ( input wire [31:0] x,
      output reg [31:0] y,
      input wire clk,
      input wire rstn
);

    wire s;
    wire [7:0] e;
    wire [22:0] m;
    wire [35:0] val;
    wire [9:0] key;
    wire [31:0] y_wire;

    reg reg_s;
    reg [7:0] reg_e;
    reg [22:0] reg_m;
    reg [22:0] reg_c;
    reg [12:0] reg_d;

    assign s = x[31];
    assign e = x[30:23];
    assign m = x[22:0];
    assign key = m[22:13];

    finv_table u1(key, val, clk, rstn);
    finv_1st u2(reg_s, reg_e, reg_m, reg_c, reg_d, y_wire);

    always @(posedge clk) begin
        reg_c <= val[35:13];
        reg_d <= val[12:0];
        reg_s <= s;
        reg_e <= e;
        reg_m <= m;
        y <= y_wire;
    end

endmodule


module finv_1st
    (input wire s,
     input wire [7:0] e,
     input wire [22:0] m,
     input wire [22:0] c,
     input wire [12:0] d,
     output wire [31:0] y);

    wire f;
    wire [9:0] a0;
    wire [12:0] a1;
    wire [25:0] cor_n;
    wire [13:0] cor;
    wire [22:0] ans_m;
    wire [7:0] e0;
    wire [7:0] e1;
    wire [7:0] ans_e;

    assign a0 = m[22:13];
    assign a1 = m[12:0];
    assign cor_n = a1 * d;
    assign cor = (a0 < 10'd424) ? (cor_n >> 12) : (cor_n >> 13);
    assign ans_m = c - cor;
    assign f = (m == 23'b0) ? 0 : 1;
    assign e0 = 8'd254 - e;
    assign e1 = e0 - f;
    assign ans_e = (e == 0) ? 0 : e1;
    assign y = {s, ans_e, ans_m};

endmodule


module finv_table
    (input wire [9:0] addr,
     output reg [35:0] dout,
     input wire clk,
     input wire rstn
);

    reg [35:0] finv_table [1023:0];

initial
    begin
        finv_table[1023] = 36'h002003001;
        finv_table[1022] = 36'h00400F006;
        finv_table[1021] = 36'h00602300A;
        finv_table[1020] = 36'h00803F00E;
        finv_table[1019] = 36'h00A063012;
        finv_table[1018] = 36'h00C08F015;
        finv_table[1017] = 36'h00E0C3019;
        finv_table[1016] = 36'h0100FF01D;
        finv_table[1015] = 36'h012143022;
        finv_table[1014] = 36'h01418F026;
        finv_table[1013] = 36'h0161E502B;
        finv_table[1012] = 36'h01824102D;
        finv_table[1011] = 36'h01A2A7032;
        finv_table[1010] = 36'h01C313035;
        finv_table[1009] = 36'h01E38903A;
        finv_table[1008] = 36'h02040703E;
        finv_table[1007] = 36'h02248B041;
        finv_table[1006] = 36'h024519047;
        finv_table[1005] = 36'h0265AF04B;
        finv_table[1004] = 36'h02864D04F;
        finv_table[1003] = 36'h02A6F5053;
        finv_table[1002] = 36'h02C7A3056;
        finv_table[1001] = 36'h02E85B05B;
        finv_table[1000] = 36'h030919060;
        finv_table[999] = 36'h0329E1064;
        finv_table[998] = 36'h034AB1067;
        finv_table[997] = 36'h036B8906B;
        finv_table[996] = 36'h038C69070;
        finv_table[995] = 36'h03AD53074;
        finv_table[994] = 36'h03CE43077;
        finv_table[993] = 36'h03EF3D07D;
        finv_table[992] = 36'h04103F081;
        finv_table[991] = 36'h043149085;
        finv_table[990] = 36'h04525D089;
        finv_table[989] = 36'h04737708E;
        finv_table[988] = 36'h04949B091;
        finv_table[987] = 36'h04B5C7095;
        finv_table[986] = 36'h04D6FB099;
        finv_table[985] = 36'h04F83909E;
        finv_table[984] = 36'h05197D0A1;
        finv_table[983] = 36'h053ACB0A7;
        finv_table[982] = 36'h055C210AB;
        finv_table[981] = 36'h057D810B0;
        finv_table[980] = 36'h059EE90B3;
        finv_table[979] = 36'h05C0570B8;
        finv_table[978] = 36'h05E1D10BD;
        finv_table[977] = 36'h0603510BF;
        finv_table[976] = 36'h0624DB0C5;
        finv_table[975] = 36'h06466D0C9;
        finv_table[974] = 36'h0668090CD;
        finv_table[973] = 36'h0689AB0D0;
        finv_table[972] = 36'h06AB570D6;
        finv_table[971] = 36'h06CD0D0DA;
        finv_table[970] = 36'h06EEC90DE;
        finv_table[969] = 36'h07108F0E3;
        finv_table[968] = 36'h07325F0E8;
        finv_table[967] = 36'h0754370EB;
        finv_table[966] = 36'h0776170F0;
        finv_table[965] = 36'h0797FF0F3;
        finv_table[964] = 36'h07B9F10F8;
        finv_table[963] = 36'h07DBEB0FC;
        finv_table[962] = 36'h07FDEF101;
        finv_table[961] = 36'h081FF9106;
        finv_table[960] = 36'h08420F10A;
        finv_table[959] = 36'h08642B10E;
        finv_table[958] = 36'h088653113;
        finv_table[957] = 36'h08A881116;
        finv_table[956] = 36'h08CAB911C;
        finv_table[955] = 36'h08ECF9120;
        finv_table[954] = 36'h090F43125;
        finv_table[953] = 36'h093197129;
        finv_table[952] = 36'h0953F112C;
        finv_table[951] = 36'h097655132;
        finv_table[950] = 36'h0998C3137;
        finv_table[949] = 36'h09BB3913B;
        finv_table[948] = 36'h09DDB913F;
        finv_table[947] = 36'h0A0041143;
        finv_table[946] = 36'h0A22D1147;
        finv_table[945] = 36'h0A456B14D;
        finv_table[944] = 36'h0A680F151;
        finv_table[943] = 36'h0A8ABB155;
        finv_table[942] = 36'h0AAD6F15A;
        finv_table[941] = 36'h0AD02D15F;
        finv_table[940] = 36'h0AF2F5164;
        finv_table[939] = 36'h0B15C5168;
        finv_table[938] = 36'h0B389F16C;
        finv_table[937] = 36'h0B5B81170;
        finv_table[936] = 36'h0B7E6D175;
        finv_table[935] = 36'h0BA161179;
        finv_table[934] = 36'h0BC45F17F;
        finv_table[933] = 36'h0BE767183;
        finv_table[932] = 36'h0C0A77188;
        finv_table[931] = 36'h0C2D8F18B;
        finv_table[930] = 36'h0C50B3191;
        finv_table[929] = 36'h0C73DF196;
        finv_table[928] = 36'h0C971319B;
        finv_table[927] = 36'h0CBA5119E;
        finv_table[926] = 36'h0CDD991A3;
        finv_table[925] = 36'h0D00E91A7;
        finv_table[924] = 36'h0D24431AD;
        finv_table[923] = 36'h0D47A71B1;
        finv_table[922] = 36'h0D6B131B5;
        finv_table[921] = 36'h0D8E891BB;
        finv_table[920] = 36'h0DB2091BF;
        finv_table[919] = 36'h0DD5911C3;
        finv_table[918] = 36'h0DF9231C9;
        finv_table[917] = 36'h0E1CBF1CD;
        finv_table[916] = 36'h0E40631D1;
        finv_table[915] = 36'h0E64111D7;
        finv_table[914] = 36'h0E87C91DC;
        finv_table[913] = 36'h0EAB8B1E0;
        finv_table[912] = 36'h0ECF551E5;
        finv_table[911] = 36'h0EF3291E9;
        finv_table[910] = 36'h0F17071EE;
        finv_table[909] = 36'h0F3AED1F2;
        finv_table[908] = 36'h0F5EDD1F8;
        finv_table[907] = 36'h0F82D71FD;
        finv_table[906] = 36'h0FA6DB202;
        finv_table[905] = 36'h0FCAE9206;
        finv_table[904] = 36'h0FEEFF20A;
        finv_table[903] = 36'h10131F210;
        finv_table[902] = 36'h103749215;
        finv_table[901] = 36'h105B7D219;
        finv_table[900] = 36'h107FB921E;
        finv_table[899] = 36'h10A401223;
        finv_table[898] = 36'h10C851227;
        finv_table[897] = 36'h10ECAB22C;
        finv_table[896] = 36'h11110F231;
        finv_table[895] = 36'h11357D236;
        finv_table[894] = 36'h1159F323A;
        finv_table[893] = 36'h117E75241;
        finv_table[892] = 36'h11A2FF244;
        finv_table[891] = 36'h11C79524A;
        finv_table[890] = 36'h11EC3324F;
        finv_table[889] = 36'h1210DB253;
        finv_table[888] = 36'h12358D258;
        finv_table[887] = 36'h125A4925E;
        finv_table[886] = 36'h127F0D261;
        finv_table[885] = 36'h12A3DD268;
        finv_table[884] = 36'h12C8B726C;
        finv_table[883] = 36'h12ED99270;
        finv_table[882] = 36'h131287277;
        finv_table[881] = 36'h13377F27B;
        finv_table[880] = 36'h135C7F280;
        finv_table[879] = 36'h13818B285;
        finv_table[878] = 36'h13A69F28B;
        finv_table[877] = 36'h13CBBD28F;
        finv_table[876] = 36'h13F0E7295;
        finv_table[875] = 36'h141619299;
        finv_table[874] = 36'h143B5729E;
        finv_table[873] = 36'h14609D2A2;
        finv_table[872] = 36'h1485EF2A9;
        finv_table[871] = 36'h14AB4B2AD;
        finv_table[870] = 36'h14D0AF2B3;
        finv_table[869] = 36'h14F61F2B7;
        finv_table[868] = 36'h151B992BC;
        finv_table[867] = 36'h15411B2C0;
        finv_table[866] = 36'h1566A92C7;
        finv_table[865] = 36'h158C412CC;
        finv_table[864] = 36'h15B1E32D1;
        finv_table[863] = 36'h15D7912D6;
        finv_table[862] = 36'h15FD472DA;
        finv_table[861] = 36'h1623072E0;
        finv_table[860] = 36'h1648D32E6;
        finv_table[859] = 36'h166EA92EA;
        finv_table[858] = 36'h1694892F0;
        finv_table[857] = 36'h16BA732F5;
        finv_table[856] = 36'h16E0672FA;
        finv_table[855] = 36'h1706652FE;
        finv_table[854] = 36'h172C6F304;
        finv_table[853] = 36'h175281308;
        finv_table[852] = 36'h17789F30F;
        finv_table[851] = 36'h179EC7314;
        finv_table[850] = 36'h17C4FB319;
        finv_table[849] = 36'h17EB3731D;
        finv_table[848] = 36'h18117F324;
        finv_table[847] = 36'h1837D1328;
        finv_table[846] = 36'h185E2D32E;
        finv_table[845] = 36'h188495333;
        finv_table[844] = 36'h18AB07338;
        finv_table[843] = 36'h18D18333E;
        finv_table[842] = 36'h18F809343;
        finv_table[841] = 36'h191E9B348;
        finv_table[840] = 36'h19453734E;
        finv_table[839] = 36'h196BDD353;
        finv_table[838] = 36'h19928D357;
        finv_table[837] = 36'h19B94935E;
        finv_table[836] = 36'h19E00F363;
        finv_table[835] = 36'h1A06E1368;
        finv_table[834] = 36'h1A2DBD36D;
        finv_table[833] = 36'h1A54A3372;
        finv_table[832] = 36'h1A7B95378;
        finv_table[831] = 36'h1AA29137E;
        finv_table[830] = 36'h1AC997383;
        finv_table[829] = 36'h1AF0A9388;
        finv_table[828] = 36'h1B17C538E;
        finv_table[827] = 36'h1B3EEB392;
        finv_table[826] = 36'h1B661D399;
        finv_table[825] = 36'h1B8D5B39E;
        finv_table[824] = 36'h1BB4A33A4;
        finv_table[823] = 36'h1BDBF53A9;
        finv_table[822] = 36'h1C03533AF;
        finv_table[821] = 36'h1C2ABB3B4;
        finv_table[820] = 36'h1C522D3B8;
        finv_table[819] = 36'h1C79AD3BF;
        finv_table[818] = 36'h1CA1353C5;
        finv_table[817] = 36'h1CC8C93CA;
        finv_table[816] = 36'h1CF0693CF;
        finv_table[815] = 36'h1D18133D4;
        finv_table[814] = 36'h1D3FC93DA;
        finv_table[813] = 36'h1D67893DF;
        finv_table[812] = 36'h1D8F553E5;
        finv_table[811] = 36'h1DB72B3EA;
        finv_table[810] = 36'h1DDF0D3F0;
        finv_table[809] = 36'h1E06F93F5;
        finv_table[808] = 36'h1E2EF13FC;
        finv_table[807] = 36'h1E56F5401;
        finv_table[806] = 36'h1E7F03406;
        finv_table[805] = 36'h1EA71D40C;
        finv_table[804] = 36'h1ECF41411;
        finv_table[803] = 36'h1EF771418;
        finv_table[802] = 36'h1F1FAD41E;
        finv_table[801] = 36'h1F47F3423;
        finv_table[800] = 36'h1F7045429;
        finv_table[799] = 36'h1F98A342F;
        finv_table[798] = 36'h1FC10B434;
        finv_table[797] = 36'h1FE97F43A;
        finv_table[796] = 36'h2011FF440;
        finv_table[795] = 36'h203A89445;
        finv_table[794] = 36'h20632144B;
        finv_table[793] = 36'h208BC1450;
        finv_table[792] = 36'h20B46F456;
        finv_table[791] = 36'h20DD2745B;
        finv_table[790] = 36'h2105EB461;
        finv_table[789] = 36'h212EBB467;
        finv_table[788] = 36'h21579746E;
        finv_table[787] = 36'h21807D473;
        finv_table[786] = 36'h21A96F478;
        finv_table[785] = 36'h21D26D47E;
        finv_table[784] = 36'h21FB77485;
        finv_table[783] = 36'h22248B48A;
        finv_table[782] = 36'h224DAB48F;
        finv_table[781] = 36'h2276D9496;
        finv_table[780] = 36'h22A01149C;
        finv_table[779] = 36'h22C9534A1;
        finv_table[778] = 36'h22F2A34A8;
        finv_table[777] = 36'h231BFF4AD;
        finv_table[776] = 36'h2345654B2;
        finv_table[775] = 36'h236ED94B9;
        finv_table[774] = 36'h2398574BF;
        finv_table[773] = 36'h23C1E14C4;
        finv_table[772] = 36'h23EB774CA;
        finv_table[771] = 36'h2415194D1;
        finv_table[770] = 36'h243EC74D7;
        finv_table[769] = 36'h2468814DC;
        finv_table[768] = 36'h2492474E2;
        finv_table[767] = 36'h24BC194E8;
        finv_table[766] = 36'h24E5F74EE;
        finv_table[765] = 36'h250FE14F5;
        finv_table[764] = 36'h2539D54F9;
        finv_table[763] = 36'h2563D7501;
        finv_table[762] = 36'h258DE5506;
        finv_table[761] = 36'h25B7FF50C;
        finv_table[760] = 36'h25E225512;
        finv_table[759] = 36'h260C57518;
        finv_table[758] = 36'h26369551E;
        finv_table[757] = 36'h2660DF524;
        finv_table[756] = 36'h268B3552B;
        finv_table[755] = 36'h26B599531;
        finv_table[754] = 36'h26E007537;
        finv_table[753] = 36'h270A8353D;
        finv_table[752] = 36'h273509543;
        finv_table[751] = 36'h275F9D549;
        finv_table[750] = 36'h278A3D54F;
        finv_table[749] = 36'h27B4E9555;
        finv_table[748] = 36'h27DFA155B;
        finv_table[747] = 36'h280A67562;
        finv_table[746] = 36'h283537567;
        finv_table[745] = 36'h28601556E;
        finv_table[744] = 36'h288AFF574;
        finv_table[743] = 36'h28B5F557A;
        finv_table[742] = 36'h28E0F9581;
        finv_table[741] = 36'h290C07586;
        finv_table[740] = 36'h29372358E;
        finv_table[739] = 36'h29624D594;
        finv_table[738] = 36'h298D8159A;
        finv_table[737] = 36'h29B8C35A0;
        finv_table[736] = 36'h29E4115A7;
        finv_table[735] = 36'h2A0F6B5AC;
        finv_table[734] = 36'h2A3AD35B3;
        finv_table[733] = 36'h2A66475BA;
        finv_table[732] = 36'h2A91C75BF;
        finv_table[731] = 36'h2ABD555C6;
        finv_table[730] = 36'h2AE8EF5CD;
        finv_table[729] = 36'h2B14955D2;
        finv_table[728] = 36'h2B40495D9;
        finv_table[727] = 36'h2B6C095DF;
        finv_table[726] = 36'h2B97D75E6;
        finv_table[725] = 36'h2BC3B15ED;
        finv_table[724] = 36'h2BEF975F3;
        finv_table[723] = 36'h2C1B8B5F9;
        finv_table[722] = 36'h2C478B600;
        finv_table[721] = 36'h2C7399606;
        finv_table[720] = 36'h2C9FB360D;
        finv_table[719] = 36'h2CCBDB614;
        finv_table[718] = 36'h2CF80F61A;
        finv_table[717] = 36'h2D244F61F;
        finv_table[716] = 36'h2D509F627;
        finv_table[715] = 36'h2D7CF962E;
        finv_table[714] = 36'h2DA961634;
        finv_table[713] = 36'h2DD5D763A;
        finv_table[712] = 36'h2E025B641;
        finv_table[711] = 36'h2E2EE9648;
        finv_table[710] = 36'h2E5B8764E;
        finv_table[709] = 36'h2E8831655;
        finv_table[708] = 36'h2EB4E965C;
        finv_table[707] = 36'h2EE1AD662;
        finv_table[706] = 36'h2F0E7F669;
        finv_table[705] = 36'h2F3B5D66F;
        finv_table[704] = 36'h2F6849676;
        finv_table[703] = 36'h2F954367D;
        finv_table[702] = 36'h2FC24B683;
        finv_table[701] = 36'h2FEF5F68A;
        finv_table[700] = 36'h301C81690;
        finv_table[699] = 36'h3049AF696;
        finv_table[698] = 36'h3076ED69E;
        finv_table[697] = 36'h30A4376A5;
        finv_table[696] = 36'h30D18F6AC;
        finv_table[695] = 36'h30FEF36B2;
        finv_table[694] = 36'h312C656B8;
        finv_table[693] = 36'h3159E56C0;
        finv_table[692] = 36'h3187736C7;
        finv_table[691] = 36'h31B50F6CD;
        finv_table[690] = 36'h31E2B76D3;
        finv_table[689] = 36'h32106F6DB;
        finv_table[688] = 36'h323E336E2;
        finv_table[687] = 36'h326C056E9;
        finv_table[686] = 36'h3299E56F0;
        finv_table[685] = 36'h32C7D16F6;
        finv_table[684] = 36'h32F5CD6FD;
        finv_table[683] = 36'h3323D5703;
        finv_table[682] = 36'h3351ED70B;
        finv_table[681] = 36'h338011712;
        finv_table[680] = 36'h33AE43718;
        finv_table[679] = 36'h33DC85720;
        finv_table[678] = 36'h340AD3727;
        finv_table[677] = 36'h34392F72E;
        finv_table[676] = 36'h346799735;
        finv_table[675] = 36'h34961173C;
        finv_table[674] = 36'h34C497742;
        finv_table[673] = 36'h34F32B749;
        finv_table[672] = 36'h3521CD750;
        finv_table[671] = 36'h35507F758;
        finv_table[670] = 36'h357F3D75F;
        finv_table[669] = 36'h35AE09766;
        finv_table[668] = 36'h35DCE376C;
        finv_table[667] = 36'h360BCD774;
        finv_table[666] = 36'h363AC577C;
        finv_table[665] = 36'h3669C9782;
        finv_table[664] = 36'h3698DD789;
        finv_table[663] = 36'h36C7FF790;
        finv_table[662] = 36'h36F72F797;
        finv_table[661] = 36'h37266F79F;
        finv_table[660] = 36'h3755BB7A6;
        finv_table[659] = 36'h3785177AE;
        finv_table[658] = 36'h37B4817B5;
        finv_table[657] = 36'h37E3F97BC;
        finv_table[656] = 36'h38137F7C3;
        finv_table[655] = 36'h3843157CB;
        finv_table[654] = 36'h3872B97D2;
        finv_table[653] = 36'h38A26B7D9;
        finv_table[652] = 36'h38D22B7E0;
        finv_table[651] = 36'h3901FB7E7;
        finv_table[650] = 36'h3931D97EF;
        finv_table[649] = 36'h3961C57F6;
        finv_table[648] = 36'h3991C17FD;
        finv_table[647] = 36'h39C1CB805;
        finv_table[646] = 36'h39F1E380B;
        finv_table[645] = 36'h3A220B813;
        finv_table[644] = 36'h3A524181A;
        finv_table[643] = 36'h3A8287822;
        finv_table[642] = 36'h3AB2DB82A;
        finv_table[641] = 36'h3AE33D831;
        finv_table[640] = 36'h3B13AF838;
        finv_table[639] = 36'h3B442F83F;
        finv_table[638] = 36'h3B74BF847;
        finv_table[637] = 36'h3BA55F850;
        finv_table[636] = 36'h3BD60B856;
        finv_table[635] = 36'h3C06C985F;
        finv_table[634] = 36'h3C3793865;
        finv_table[633] = 36'h3C686F86D;
        finv_table[632] = 36'h3C9959875;
        finv_table[631] = 36'h3CCA5187C;
        finv_table[630] = 36'h3CFB59883;
        finv_table[629] = 36'h3D2C7188B;
        finv_table[628] = 36'h3D5D97893;
        finv_table[627] = 36'h3D8ECD89B;
        finv_table[626] = 36'h3DC0118A1;
        finv_table[625] = 36'h3DF1678AA;
        finv_table[624] = 36'h3E22C98B1;
        finv_table[623] = 36'h3E543D8B9;
        finv_table[622] = 36'h3E85BF8C1;
        finv_table[621] = 36'h3EB7518C8;
        finv_table[620] = 36'h3EE8F38D1;
        finv_table[619] = 36'h3F1AA38D8;
        finv_table[618] = 36'h3F4C638E0;
        finv_table[617] = 36'h3F7E338E8;
        finv_table[616] = 36'h3FB0118EE;
        finv_table[615] = 36'h3FE2018F7;
        finv_table[614] = 36'h4013FF8FF;
        finv_table[613] = 36'h40460D906;
        finv_table[612] = 36'h40782B90E;
        finv_table[611] = 36'h40AA59917;
        finv_table[610] = 36'h40DC9591E;
        finv_table[609] = 36'h410EE3926;
        finv_table[608] = 36'h41413F92E;
        finv_table[607] = 36'h4173AB935;
        finv_table[606] = 36'h41A62993F;
        finv_table[605] = 36'h41D8B5946;
        finv_table[604] = 36'h420B5194E;
        finv_table[603] = 36'h423DFD956;
        finv_table[602] = 36'h4270B995E;
        finv_table[601] = 36'h42A385966;
        finv_table[600] = 36'h42D66196E;
        finv_table[599] = 36'h43094D976;
        finv_table[598] = 36'h433C4997E;
        finv_table[597] = 36'h436F55986;
        finv_table[596] = 36'h43A27198E;
        finv_table[595] = 36'h43D59D995;
        finv_table[594] = 36'h4408DB99F;
        finv_table[593] = 36'h443C279A6;
        finv_table[592] = 36'h446F859AF;
        finv_table[591] = 36'h44A2F19B6;
        finv_table[590] = 36'h44D66F9BE;
        finv_table[589] = 36'h4509FD9C6;
        finv_table[588] = 36'h453D9D9D0;
        finv_table[587] = 36'h45714B9D7;
        finv_table[586] = 36'h45A50B9E0;
        finv_table[585] = 36'h45D8DB9E8;
        finv_table[584] = 36'h460CBB9F0;
        finv_table[583] = 36'h4640AB9F8;
        finv_table[582] = 36'h4674ADA00;
        finv_table[581] = 36'h46A8BFA09;
        finv_table[580] = 36'h46DCE1A11;
        finv_table[579] = 36'h471115A1A;
        finv_table[578] = 36'h474559A22;
        finv_table[577] = 36'h4779ADA2A;
        finv_table[576] = 36'h47AE13A33;
        finv_table[575] = 36'h47E289A3B;
        finv_table[574] = 36'h48170FA43;
        finv_table[573] = 36'h484BA7A4B;
        finv_table[572] = 36'h488051A55;
        finv_table[571] = 36'h48B509A5C;
        finv_table[570] = 36'h48E9D5A66;
        finv_table[569] = 36'h491EAFA6D;
        finv_table[568] = 36'h49539DA77;
        finv_table[567] = 36'h498899A7E;
        finv_table[566] = 36'h49BDA9A88;
        finv_table[565] = 36'h49F2C9A90;
        finv_table[564] = 36'h4A27F9A98;
        finv_table[563] = 36'h4A5D3BAA1;
        finv_table[562] = 36'h4A928DAA9;
        finv_table[561] = 36'h4AC7F3AB2;
        finv_table[560] = 36'h4AFD69ABB;
        finv_table[559] = 36'h4B32EFAC3;
        finv_table[558] = 36'h4B6887ACC;
        finv_table[557] = 36'h4B9E31AD5;
        finv_table[556] = 36'h4BD3EBADD;
        finv_table[555] = 36'h4C09B9AE7;
        finv_table[554] = 36'h4C3F97AEF;
        finv_table[553] = 36'h4C7585AF7;
        finv_table[552] = 36'h4CAB87B01;
        finv_table[551] = 36'h4CE199B09;
        finv_table[550] = 36'h4D17BDB12;
        finv_table[549] = 36'h4D4DF3B1B;
        finv_table[548] = 36'h4D8439B23;
        finv_table[547] = 36'h4DBA93B2C;
        finv_table[546] = 36'h4DF0FDB35;
        finv_table[545] = 36'h4E277BB3F;
        finv_table[544] = 36'h4E5E09B47;
        finv_table[543] = 36'h4E94A9B50;
        finv_table[542] = 36'h4ECB5BB59;
        finv_table[541] = 36'h4F021FB62;
        finv_table[540] = 36'h4F38F5B6B;
        finv_table[539] = 36'h4F6FDBB73;
        finv_table[538] = 36'h4FA6D5B7C;
        finv_table[537] = 36'h4FDDE1B85;
        finv_table[536] = 36'h5014FFB8E;
        finv_table[535] = 36'h504C2FB98;
        finv_table[534] = 36'h508371BA1;
        finv_table[533] = 36'h50BAC5BA9;
        finv_table[532] = 36'h50F22DBB4;
        finv_table[531] = 36'h5129A5BBC;
        finv_table[530] = 36'h51612FBC5;
        finv_table[529] = 36'h5198CDBCE;
        finv_table[528] = 36'h51D07DBD8;
        finv_table[527] = 36'h52083FBE1;
        finv_table[526] = 36'h524013BEA;
        finv_table[525] = 36'h5277FBBF4;
        finv_table[524] = 36'h52AFF3BFC;
        finv_table[523] = 36'h52E7FFC06;
        finv_table[522] = 36'h53201DC0E;
        finv_table[521] = 36'h53584FC19;
        finv_table[520] = 36'h539093C22;
        finv_table[519] = 36'h53C8E9C2B;
        finv_table[518] = 36'h540153C35;
        finv_table[517] = 36'h5439CDC3D;
        finv_table[516] = 36'h54725DC48;
        finv_table[515] = 36'h54AAFDC50;
        finv_table[514] = 36'h54E3B3C5B;
        finv_table[513] = 36'h551C79C63;
        finv_table[512] = 36'h555553C6D;
        finv_table[511] = 36'h558E41C77;
        finv_table[510] = 36'h55C741C80;
        finv_table[509] = 36'h560053C89;
        finv_table[508] = 36'h563979C92;
        finv_table[507] = 36'h5672B3C9D;
        finv_table[506] = 36'h56ABFFCA6;
        finv_table[505] = 36'h56E55FCB0;
        finv_table[504] = 36'h571ED1CB9;
        finv_table[503] = 36'h575857CC2;
        finv_table[502] = 36'h5791F1CCC;
        finv_table[501] = 36'h57CB9DCD5;
        finv_table[500] = 36'h58055FCE1;
        finv_table[499] = 36'h583F31CE9;
        finv_table[498] = 36'h587919CF4;
        finv_table[497] = 36'h58B313CFD;
        finv_table[496] = 36'h58ED21D07;
        finv_table[495] = 36'h592743D11;
        finv_table[494] = 36'h596177D1A;
        finv_table[493] = 36'h599BC1D25;
        finv_table[492] = 36'h59D61DD2E;
        finv_table[491] = 36'h5A108DD38;
        finv_table[490] = 36'h5A4B11D42;
        finv_table[489] = 36'h5A85A9D4C;
        finv_table[488] = 36'h5AC055D56;
        finv_table[487] = 36'h5AFB13D5F;
        finv_table[486] = 36'h5B35E7D69;
        finv_table[485] = 36'h5B70CFD74;
        finv_table[484] = 36'h5BABCBD7E;
        finv_table[483] = 36'h5BE6D9D87;
        finv_table[482] = 36'h5C21FDD91;
        finv_table[481] = 36'h5C5D35D9C;
        finv_table[480] = 36'h5C9881DA6;
        finv_table[479] = 36'h5CD3E1DB0;
        finv_table[478] = 36'h5D0F55DBA;
        finv_table[477] = 36'h5D4ADDDC4;
        finv_table[476] = 36'h5D867BDCF;
        finv_table[475] = 36'h5DC22BDD8;
        finv_table[474] = 36'h5DFDF1DE3;
        finv_table[473] = 36'h5E39CBDED;
        finv_table[472] = 36'h5E75B9DF7;
        finv_table[471] = 36'h5EB1BDE02;
        finv_table[470] = 36'h5EEDD3E0B;
        finv_table[469] = 36'h5F29FFE15;
        finv_table[468] = 36'h5F6641E20;
        finv_table[467] = 36'h5FA297E2B;
        finv_table[466] = 36'h5FDF01E35;
        finv_table[465] = 36'h601B81E40;
        finv_table[464] = 36'h605813E49;
        finv_table[463] = 36'h6094BDE55;
        finv_table[462] = 36'h60D179E5E;
        finv_table[461] = 36'h610E4DE69;
        finv_table[460] = 36'h614B35E74;
        finv_table[459] = 36'h618831E7E;
        finv_table[458] = 36'h61C543E89;
        finv_table[457] = 36'h620269E93;
        finv_table[456] = 36'h623FA5E9E;
        finv_table[455] = 36'h627CF7EA9;
        finv_table[454] = 36'h62BA5DEB3;
        finv_table[453] = 36'h62F7D9EBE;
        finv_table[452] = 36'h633569EC8;
        finv_table[451] = 36'h63730FED3;
        finv_table[450] = 36'h63B0CBEDD;
        finv_table[449] = 36'h63EE9DEE9;
        finv_table[448] = 36'h642C83EF3;
        finv_table[447] = 36'h646A7FEFE;
        finv_table[446] = 36'h64A891F09;
        finv_table[445] = 36'h64E6B9F14;
        finv_table[444] = 36'h6524F7F1F;
        finv_table[443] = 36'h656349F29;
        finv_table[442] = 36'h65A1B1F34;
        finv_table[441] = 36'h65E031F40;
        finv_table[440] = 36'h661EC3F49;
        finv_table[439] = 36'h665D6FF55;
        finv_table[438] = 36'h669C2FF60;
        finv_table[437] = 36'h66DB05F6B;
        finv_table[436] = 36'h6719F1F76;
        finv_table[435] = 36'h6758F3F81;
        finv_table[434] = 36'h67980DF8D;
        finv_table[433] = 36'h67D739F96;
        finv_table[432] = 36'h68167FFA2;
        finv_table[431] = 36'h6855DBFAE;
        finv_table[430] = 36'h68954BFB8;
        finv_table[429] = 36'h68D4D3FC4;
        finv_table[428] = 36'h691471FCF;
        finv_table[427] = 36'h695427FDB;
        finv_table[426] = 36'h6993EFFE4;
        finv_table[425] = 36'h69D3D3FF1;
        finv_table[424] = 36'h6A13CBFFC;
        finv_table[423] = 36'h6A53D9004;
        finv_table[422] = 36'h6A93FD009;
        finv_table[421] = 36'h6AD43B00F;
        finv_table[420] = 36'h6B148F015;
        finv_table[419] = 36'h6B54F701A;
        finv_table[418] = 36'h6B9577020;
        finv_table[417] = 36'h6BD611026;
        finv_table[416] = 36'h6C16BD02B;
        finv_table[415] = 36'h6C5783031;
        finv_table[414] = 36'h6C9861037;
        finv_table[413] = 36'h6CD95503D;
        finv_table[412] = 36'h6D1A61043;
        finv_table[411] = 36'h6D5B81048;
        finv_table[410] = 36'h6D9CBB04E;
        finv_table[409] = 36'h6DDE0B054;
        finv_table[408] = 36'h6E1F7305A;
        finv_table[407] = 36'h6E60F3060;
        finv_table[406] = 36'h6EA289065;
        finv_table[405] = 36'h6EE43706B;
        finv_table[404] = 36'h6F25FD071;
        finv_table[403] = 36'h6F67DB077;
        finv_table[402] = 36'h6FA9D107D;
        finv_table[401] = 36'h6FEBDD083;
        finv_table[400] = 36'h702E03089;
        finv_table[399] = 36'h70703F08F;
        finv_table[398] = 36'h70B293095;
        finv_table[397] = 36'h70F4FF09B;
        finv_table[396] = 36'h7137830A1;
        finv_table[395] = 36'h717A1F0A7;
        finv_table[394] = 36'h71BCD50AD;
        finv_table[393] = 36'h71FFA10B3;
        finv_table[392] = 36'h7242850B9;
        finv_table[391] = 36'h7285810BF;
        finv_table[390] = 36'h72C8970C5;
        finv_table[389] = 36'h730BC30CB;
        finv_table[388] = 36'h734F090D1;
        finv_table[387] = 36'h7392670D7;
        finv_table[386] = 36'h73D5DD0DD;
        finv_table[385] = 36'h74196B0E3;
        finv_table[384] = 36'h745D150EA;
        finv_table[383] = 36'h74A0D50F0;
        finv_table[382] = 36'h74E4AD0F6;
        finv_table[381] = 36'h75289D0FC;
        finv_table[380] = 36'h756CA9103;
        finv_table[379] = 36'h75B0CB108;
        finv_table[378] = 36'h75F50910F;
        finv_table[377] = 36'h76395D115;
        finv_table[376] = 36'h767DCB11B;
        finv_table[375] = 36'h76C251121;
        finv_table[374] = 36'h7706F3128;
        finv_table[373] = 36'h774BAB12E;
        finv_table[372] = 36'h77907D134;
        finv_table[371] = 36'h77D56913B;
        finv_table[370] = 36'h781A6F141;
        finv_table[369] = 36'h785F8D148;
        finv_table[368] = 36'h78A4C514E;
        finv_table[367] = 36'h78EA15154;
        finv_table[366] = 36'h792F8115B;
        finv_table[365] = 36'h797505161;
        finv_table[364] = 36'h79BAA3167;
        finv_table[363] = 36'h7A005B16E;
        finv_table[362] = 36'h7A462D174;
        finv_table[361] = 36'h7A8C1917B;
        finv_table[360] = 36'h7AD21D181;
        finv_table[359] = 36'h7B183B187;
        finv_table[358] = 36'h7B5E7518E;
        finv_table[357] = 36'h7BA4C7194;
        finv_table[356] = 36'h7BEB3519B;
        finv_table[355] = 36'h7C31BD1A2;
        finv_table[354] = 36'h7C785F1A8;
        finv_table[353] = 36'h7CBF191AE;
        finv_table[352] = 36'h7D05F11B6;
        finv_table[351] = 36'h7D4CE11BC;
        finv_table[350] = 36'h7D93EB1C2;
        finv_table[349] = 36'h7DDB111C9;
        finv_table[348] = 36'h7E22511D0;
        finv_table[347] = 36'h7E69AB1D6;
        finv_table[346] = 36'h7EB1211DD;
        finv_table[345] = 36'h7EF8B11E4;
        finv_table[344] = 36'h7F405B1EA;
        finv_table[343] = 36'h7F88211F1;
        finv_table[342] = 36'h7FD0031F8;
        finv_table[341] = 36'h8017FF1FF;
        finv_table[340] = 36'h806015206;
        finv_table[339] = 36'h80A84520C;
        finv_table[338] = 36'h80F093213;
        finv_table[337] = 36'h8138FB21A;
        finv_table[336] = 36'h81817D220;
        finv_table[335] = 36'h81CA1D228;
        finv_table[334] = 36'h8212D522E;
        finv_table[333] = 36'h825BAB235;
        finv_table[332] = 36'h82A49D23C;
        finv_table[331] = 36'h82EDA9243;
        finv_table[330] = 36'h8336D124A;
        finv_table[329] = 36'h838015251;
        finv_table[328] = 36'h83C973257;
        finv_table[327] = 36'h8412EF25F;
        finv_table[326] = 36'h845C87266;
        finv_table[325] = 36'h84A63B26D;
        finv_table[324] = 36'h84F009274;
        finv_table[323] = 36'h8539F327A;
        finv_table[322] = 36'h8583FB282;
        finv_table[321] = 36'h85CE1D288;
        finv_table[320] = 36'h86185F290;
        finv_table[319] = 36'h8662B9297;
        finv_table[318] = 36'h86AD3329E;
        finv_table[317] = 36'h86F7C72A5;
        finv_table[316] = 36'h8742772AC;
        finv_table[315] = 36'h878D452B3;
        finv_table[314] = 36'h87D8312BB;
        finv_table[313] = 36'h8823392C2;
        finv_table[312] = 36'h886E5B2C9;
        finv_table[311] = 36'h88B99B2D0;
        finv_table[310] = 36'h8904F92D7;
        finv_table[309] = 36'h8950732DE;
        finv_table[308] = 36'h899C0B2E6;
        finv_table[307] = 36'h89E7C12ED;
        finv_table[306] = 36'h8A33912F4;
        finv_table[305] = 36'h8A7F812FC;
        finv_table[304] = 36'h8ACB8D303;
        finv_table[303] = 36'h8B17B730A;
        finv_table[302] = 36'h8B63FD311;
        finv_table[301] = 36'h8BB063319;
        finv_table[300] = 36'h8BFCE5321;
        finv_table[299] = 36'h8C4985328;
        finv_table[298] = 36'h8C964132F;
        finv_table[297] = 36'h8CE31B336;
        finv_table[296] = 36'h8D301533E;
        finv_table[295] = 36'h8D7D2B345;
        finv_table[294] = 36'h8DCA6134D;
        finv_table[293] = 36'h8E17B3354;
        finv_table[292] = 36'h8E652335C;
        finv_table[291] = 36'h8EB2B3364;
        finv_table[290] = 36'h8F005F36B;
        finv_table[289] = 36'h8F4E2B373;
        finv_table[288] = 36'h8F9C1537A;
        finv_table[287] = 36'h8FEA1D382;
        finv_table[286] = 36'h903843389;
        finv_table[285] = 36'h908689391;
        finv_table[284] = 36'h90D4ED399;
        finv_table[283] = 36'h91236F3A0;
        finv_table[282] = 36'h9172113A8;
        finv_table[281] = 36'h91C0D13B0;
        finv_table[280] = 36'h920FB13B8;
        finv_table[279] = 36'h925EAF3BF;
        finv_table[278] = 36'h92ADCD3C7;
        finv_table[277] = 36'h92FD093CF;
        finv_table[276] = 36'h934C633D6;
        finv_table[275] = 36'h939BDF3DF;
        finv_table[274] = 36'h93EB7B3E7;
        finv_table[273] = 36'h943B333EE;
        finv_table[272] = 36'h948B0B3F6;
        finv_table[271] = 36'h94DB053FE;
        finv_table[270] = 36'h952B1D406;
        finv_table[269] = 36'h957B5540E;
        finv_table[268] = 36'h95CBAD416;
        finv_table[267] = 36'h961C2541E;
        finv_table[266] = 36'h966CBD426;
        finv_table[265] = 36'h96BD7342E;
        finv_table[264] = 36'h970E4B436;
        finv_table[263] = 36'h975F4343E;
        finv_table[262] = 36'h97B05B446;
        finv_table[261] = 36'h98019544E;
        finv_table[260] = 36'h9852ED456;
        finv_table[259] = 36'h98A46745E;
        finv_table[258] = 36'h98F5FF466;
        finv_table[257] = 36'h9947BB46F;
        finv_table[256] = 36'h999995476;
        finv_table[255] = 36'h99EB9147F;
        finv_table[254] = 36'h9A3DAF487;
        finv_table[253] = 36'h9A8FEB48F;
        finv_table[252] = 36'h9AE24B498;
        finv_table[251] = 36'h9B34CB4A0;
        finv_table[250] = 36'h9B876B4A8;
        finv_table[249] = 36'h9BDA2D4B0;
        finv_table[248] = 36'h9C2D114B9;
        finv_table[247] = 36'h9C80154C1;
        finv_table[246] = 36'h9CD33D4CA;
        finv_table[245] = 36'h9D26834D2;
        finv_table[244] = 36'h9D79ED4DA;
        finv_table[243] = 36'h9DCD794E3;
        finv_table[242] = 36'h9E21254EB;
        finv_table[241] = 36'h9E74F54F4;
        finv_table[240] = 36'h9EC8E54FC;
        finv_table[239] = 36'h9F1CF9505;
        finv_table[238] = 36'h9F712D50D;
        finv_table[237] = 36'h9FC585516;
        finv_table[236] = 36'hA019FD51E;
        finv_table[235] = 36'hA06E99527;
        finv_table[234] = 36'hA0C35752F;
        finv_table[233] = 36'hA11839538;
        finv_table[232] = 36'hA16D3B540;
        finv_table[231] = 36'hA1C261549;
        finv_table[230] = 36'hA217AB552;
        finv_table[229] = 36'hA26D1555B;
        finv_table[228] = 36'hA2C2A5564;
        finv_table[227] = 36'hA3185756C;
        finv_table[226] = 36'hA36E2B575;
        finv_table[225] = 36'hA3C42357E;
        finv_table[224] = 36'hA41A3D586;
        finv_table[223] = 36'hA4707D590;
        finv_table[222] = 36'hA4C6DF598;
        finv_table[221] = 36'hA51D635A1;
        finv_table[220] = 36'hA5740D5AA;
        finv_table[219] = 36'hA5CAD95B3;
        finv_table[218] = 36'hA621C95BC;
        finv_table[217] = 36'hA678DF5C5;
        finv_table[216] = 36'hA6D0175CE;
        finv_table[215] = 36'hA727735D7;
        finv_table[214] = 36'hA77EF35E0;
        finv_table[213] = 36'hA7D6995E9;
        finv_table[212] = 36'hA82E615F2;
        finv_table[211] = 36'hA8864F5FB;
        finv_table[210] = 36'hA8DE61604;
        finv_table[209] = 36'hA9369760D;
        finv_table[208] = 36'hA98EF3617;
        finv_table[207] = 36'hA9E771620;
        finv_table[206] = 36'hAA4017629;
        finv_table[205] = 36'hAA98E1632;
        finv_table[204] = 36'hAAF1CF63B;
        finv_table[203] = 36'hAB4AE3645;
        finv_table[202] = 36'hABA41B64E;
        finv_table[201] = 36'hABFD7B658;
        finv_table[200] = 36'hAC56FD661;
        finv_table[199] = 36'hACB0A766A;
        finv_table[198] = 36'hAD0A75673;
        finv_table[197] = 36'hAD646967D;
        finv_table[196] = 36'hADBE83686;
        finv_table[195] = 36'hAE18C3690;
        finv_table[194] = 36'hAE7329699;
        finv_table[193] = 36'hAECDB56A3;
        finv_table[192] = 36'hAF28676AC;
        finv_table[191] = 36'hAF83416B6;
        finv_table[190] = 36'hAFDE3F6C0;
        finv_table[189] = 36'hB039636C9;
        finv_table[188] = 36'hB094AF6D3;
        finv_table[187] = 36'hB0F0216DC;
        finv_table[186] = 36'hB14BB96E6;
        finv_table[185] = 36'hB1A7796F0;
        finv_table[184] = 36'hB203616FA;
        finv_table[183] = 36'hB25F6D703;
        finv_table[182] = 36'hB2BBA170D;
        finv_table[181] = 36'hB317FD717;
        finv_table[180] = 36'hB37481721;
        finv_table[179] = 36'hB3D12B72A;
        finv_table[178] = 36'hB42DFD734;
        finv_table[177] = 36'hB48AF773E;
        finv_table[176] = 36'hB4E817748;
        finv_table[175] = 36'hB54561752;
        finv_table[174] = 36'hB5A2D175C;
        finv_table[173] = 36'hB60069766;
        finv_table[172] = 36'hB65E2B770;
        finv_table[171] = 36'hB6BC1377A;
        finv_table[170] = 36'hB71A25784;
        finv_table[169] = 36'hB7785D78E;
        finv_table[168] = 36'hB7D6BF798;
        finv_table[167] = 36'hB8354B7A3;
        finv_table[166] = 36'hB893FD7AC;
        finv_table[165] = 36'hB8F2D97B7;
        finv_table[164] = 36'hB951DF7C1;
        finv_table[163] = 36'hB9B10D7CB;
        finv_table[162] = 36'hBA10637D5;
        finv_table[161] = 36'hBA6FE37E0;
        finv_table[160] = 36'hBACF8D7EA;
        finv_table[159] = 36'hBB2F617F5;
        finv_table[158] = 36'hBB8F5D7FF;
        finv_table[157] = 36'hBBEF83809;
        finv_table[156] = 36'hBC4FD3814;
        finv_table[155] = 36'hBCB04B81E;
        finv_table[154] = 36'hBD10EF829;
        finv_table[153] = 36'hBD71BD833;
        finv_table[152] = 36'hBDD2B583E;
        finv_table[151] = 36'hBE33D7848;
        finv_table[150] = 36'hBE9523853;
        finv_table[149] = 36'hBEF69985D;
        finv_table[148] = 36'hBF583B868;
        finv_table[147] = 36'hBFBA07873;
        finv_table[146] = 36'hC01BFD87D;
        finv_table[145] = 36'hC07E1F888;
        finv_table[144] = 36'hC0E06D893;
        finv_table[143] = 36'hC142E589E;
        finv_table[142] = 36'hC1A5878A8;
        finv_table[141] = 36'hC208558B3;
        finv_table[140] = 36'hC26B4F8BE;
        finv_table[139] = 36'hC2CE758C9;
        finv_table[138] = 36'hC331C78D4;
        finv_table[137] = 36'hC395438DF;
        finv_table[136] = 36'hC3F8ED8EA;
        finv_table[135] = 36'hC45CC18F5;
        finv_table[134] = 36'hC4C0C3900;
        finv_table[133] = 36'hC524EF90B;
        finv_table[132] = 36'hC58949916;
        finv_table[131] = 36'hC5EDCF921;
        finv_table[130] = 36'hC6528192C;
        finv_table[129] = 36'hC6B761938;
        finv_table[128] = 36'hC71C6D943;
        finv_table[127] = 36'hC781A794E;
        finv_table[126] = 36'hC7E70D959;
        finv_table[125] = 36'hC84CA1965;
        finv_table[124] = 36'hC8B261970;
        finv_table[123] = 36'hC9184F97B;
        finv_table[122] = 36'hC97E6B987;
        finv_table[121] = 36'hC9E4B5992;
        finv_table[120] = 36'hCA4B2D99E;
        finv_table[119] = 36'hCAB1D19A9;
        finv_table[118] = 36'hCB18A59B5;
        finv_table[117] = 36'hCB7FA59C0;
        finv_table[116] = 36'hCBE6D59CC;
        finv_table[115] = 36'hCC4E339D7;
        finv_table[114] = 36'hCCB5BF9E3;
        finv_table[113] = 36'hCD1D7B9EF;
        finv_table[112] = 36'hCD85639FA;
        finv_table[111] = 36'hCDED7DA06;
        finv_table[110] = 36'hCE55C5A12;
        finv_table[109] = 36'hCEBE3BA1D;
        finv_table[108] = 36'hCF26E1A29;
        finv_table[107] = 36'hCF8FB7A35;
        finv_table[106] = 36'hCFF8BBA41;
        finv_table[105] = 36'hD061F1A4D;
        finv_table[104] = 36'hD0CB55A59;
        finv_table[103] = 36'hD134E9A65;
        finv_table[102] = 36'hD19EADA71;
        finv_table[101] = 36'hD208A1A7D;
        finv_table[100] = 36'hD272C5A89;
        finv_table[99] = 36'hD2DD1BA95;
        finv_table[98] = 36'hD3479FAA1;
        finv_table[97] = 36'hD3B255AAD;
        finv_table[96] = 36'hD41D3DAB9;
        finv_table[95] = 36'hD48855AC6;
        finv_table[94] = 36'hD4F39DAD2;
        finv_table[93] = 36'hD55F17ADE;
        finv_table[92] = 36'hD5CAC5AEB;
        finv_table[91] = 36'hD636A1AF7;
        finv_table[90] = 36'hD6A2ADB03;
        finv_table[89] = 36'hD70EEFB10;
        finv_table[88] = 36'hD77B61B1C;
        finv_table[87] = 36'hD7E805B29;
        finv_table[86] = 36'hD854D9B35;
        finv_table[85] = 36'hD8C1E3B42;
        finv_table[84] = 36'hD92F1FB4F;
        finv_table[83] = 36'hD99C8BB5B;
        finv_table[82] = 36'hDA0A2BB68;
        finv_table[81] = 36'hDA77FDB74;
        finv_table[80] = 36'hDAE603B81;
        finv_table[79] = 36'hDB543BB8E;
        finv_table[78] = 36'hDBC2A7B9B;
        finv_table[77] = 36'hDC3147BA8;
        finv_table[76] = 36'hDCA01BBB5;
        finv_table[75] = 36'hDD0F21BC2;
        finv_table[74] = 36'hDD7E5BBCF;
        finv_table[73] = 36'hDDEDC7BDB;
        finv_table[72] = 36'hDE5D69BE8;
        finv_table[71] = 36'hDECD3FBF5;
        finv_table[70] = 36'hDF3D4BC03;
        finv_table[69] = 36'hDFAD8BC10;
        finv_table[68] = 36'hE01DFBC1C;
        finv_table[67] = 36'hE08EA5C2A;
        finv_table[66] = 36'hE0FF83C37;
        finv_table[65] = 36'hE17097C45;
        finv_table[64] = 36'hE1E1DBC51;
        finv_table[63] = 36'hE25359C5F;
        finv_table[62] = 36'hE2C50BC6C;
        finv_table[61] = 36'hE336F5C7A;
        finv_table[60] = 36'hE3A911C87;
        finv_table[59] = 36'hE41B67C95;
        finv_table[58] = 36'hE48DEFCA2;
        finv_table[57] = 36'hE500B1CB0;
        finv_table[56] = 36'hE573A9CBE;
        finv_table[55] = 36'hE5E6D5CCB;
        finv_table[54] = 36'hE65A39CD9;
        finv_table[53] = 36'hE6CDD5CE7;
        finv_table[52] = 36'hE741A5CF4;
        finv_table[51] = 36'hE7B5ADD02;
        finv_table[50] = 36'hE829EFD10;
        finv_table[49] = 36'hE89E67D1E;
        finv_table[48] = 36'hE91317D2C;
        finv_table[47] = 36'hE987FBD39;
        finv_table[46] = 36'hE9FD1DD48;
        finv_table[45] = 36'hEA7273D56;
        finv_table[44] = 36'hEAE801D63;
        finv_table[43] = 36'hEB5DCBD72;
        finv_table[42] = 36'hEBD3CBD80;
        finv_table[41] = 36'hEC4A03D8E;
        finv_table[40] = 36'hECC075D9C;
        finv_table[39] = 36'hED3721DAB;
        finv_table[38] = 36'hEDAE05DB9;
        finv_table[37] = 36'hEE2523DC7;
        finv_table[36] = 36'hEE9C79DD5;
        finv_table[35] = 36'hEF140BDE4;
        finv_table[34] = 36'hEF8BD5DF2;
        finv_table[33] = 36'hF003DBE01;
        finv_table[32] = 36'hF07C1BE10;
        finv_table[31] = 36'hF0F493E1E;
        finv_table[30] = 36'hF16D47E2D;
        finv_table[29] = 36'hF1E635E3B;
        finv_table[28] = 36'hF25F5FE4A;
        finv_table[27] = 36'hF2D8C3E59;
        finv_table[26] = 36'hF35263E68;
        finv_table[25] = 36'hF3CC3DE76;
        finv_table[24] = 36'hF44653E85;
        finv_table[23] = 36'hF4C0A7E95;
        finv_table[22] = 36'hF53B35EA3;
        finv_table[21] = 36'hF5B5FFEB2;
        finv_table[20] = 36'hF63105EC1;
        finv_table[19] = 36'hF6AC47ED0;
        finv_table[18] = 36'hF727C7EE0;
        finv_table[17] = 36'hF7A383EEF;
        finv_table[16] = 36'hF81F7BEFE;
        finv_table[15] = 36'hF89BB3F0E;
        finv_table[14] = 36'hF91827F1D;
        finv_table[13] = 36'hF994D7F2C;
        finv_table[12] = 36'hFA11C5F3B;
        finv_table[11] = 36'hFA8EF1F4B;
        finv_table[10] = 36'hFB0C5BF5A;
        finv_table[9] = 36'hFB8A03F6A;
        finv_table[8] = 36'hFC07EBF7A;
        finv_table[7] = 36'hFC860FF89;
        finv_table[6] = 36'hFD0473F99;
        finv_table[5] = 36'hFD8317FA9;
        finv_table[4] = 36'hFE01F9FB8;
        finv_table[3] = 36'hFE8119FC8;
        finv_table[2] = 36'hFF0079FD8;
        finv_table[1] = 36'hFF8019FE8;
        finv_table[0] = 36'hFFFFFBFF8;
    end

    always @(posedge clk) begin
        dout <= finv_table[addr];
    end

endmodule

`default_nettype wire