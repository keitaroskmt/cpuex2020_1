`default_nettype none

module finv
    ( input wire [31:0] x,
      output reg [31:0] y,
      input wire clk,
      input wire rstn
);

    wire s;
    wire [7:0] e;
    wire [22:0] m;
    wire [35:0] val;
    wire [9:0] key;
    wire [31:0] y_wire;

    reg reg_s;
    reg [7:0] reg_e;
    reg [22:0] reg_m;
    reg [22:0] reg_c;
    reg [12:0] reg_d;

    assign s = x[31];
    assign e = x[30:23];
    assign m = x[22:0];
    assign key = m[22:13];

    finv_table u1(key, val, clk, rstn);
    finv_1st u2(reg_s, reg_e, reg_m, val, y_wire);

    always @(posedge clk) begin
        reg_s <= s;
        reg_e <= e;
        reg_m <= m;
        y <= y_wire;
    end

endmodule


module finv_1st
    (input wire s,
     input wire [7:0] e,
     input wire [22:0] m,
     input wire [35:0] val,
     output wire [31:0] y);

    wire [9:0] a0;
    wire [12:0] a1;
    wire [25:0] cor_n;
    wire [13:0] cor;
    wire [22:0] ans_m;
    wire [22:0] m1;
    wire [22:0] m2;
    wire [22:0] shifted_m;
    wire [7:0] e0;
    wire [7:0] e1;
    wire [7:0] ans_e;
    wire [22:0] c;
    wire [12:0] d;
    wire subnormal;
    wire [8:0] minus_e;
    wire [8:0] shift_e;

    assign c = val[35:13];
    assign d = val[12:0];
    assign a0 = m[22:13];
    assign a1 = m[12:0];
    assign cor_n = a1 * d;
    assign cor = (a0 < 10'd424) ? (cor_n >> 12) : (cor_n >> 13);
    assign e0 = 8'd254 - e;
    assign e1 = e0 - 1;
    assign minus_e = e + 1;
    assign subnormal = (e > 8'd253) ? 1 :
                       (1 >= e0) ? 1 : 0;
    assign shift_e = (subnormal == 1) ? minus_e - 254 : 0;
    assign ans_e = (e == 0) ? 0 : e1;
    assign m1 = c - cor;
    assign m2 = (m == 23'b0) ? {1'b1, 22'b0} : {1'b1, m1[22:1]};
    assign shifted_m = m2 >> shift_e;
    assign ans_m = (e == 0) ? 0 :
                   (subnormal == 1) ? shifted_m : m1;
    assign y = (subnormal == 1) ? {s, 8'b0, ans_m} : {s, ans_e, ans_m};

endmodule


module finv_table
    (input wire [9:0] addr,
     output reg [35:0] dout,
     input wire clk,
     input wire rstn
);

    reg [35:0] finv_table [1023:0];

initial
    begin
        finv_table[1023] = 36'h002003002;
        finv_table[1022] = 36'h00400F006;
        finv_table[1021] = 36'h00602300A;
        finv_table[1020] = 36'h00803F00E;
        finv_table[1019] = 36'h00A063012;
        finv_table[1018] = 36'h00C08F016;
        finv_table[1017] = 36'h00E0C301A;
        finv_table[1016] = 36'h01010101E;
        finv_table[1015] = 36'h012145023;
        finv_table[1014] = 36'h014191025;
        finv_table[1013] = 36'h0161E502A;
        finv_table[1012] = 36'h01824302E;
        finv_table[1011] = 36'h01A2A7031;
        finv_table[1010] = 36'h01C315036;
        finv_table[1009] = 36'h01E389039;
        finv_table[1008] = 36'h02040703F;
        finv_table[1007] = 36'h02248D042;
        finv_table[1006] = 36'h02451B046;
        finv_table[1005] = 36'h0265B104A;
        finv_table[1004] = 36'h02864F04E;
        finv_table[1003] = 36'h02A6F5052;
        finv_table[1002] = 36'h02C7A5057;
        finv_table[1001] = 36'h02E85B05C;
        finv_table[1000] = 36'h03091B05F;
        finv_table[999] = 36'h0329E1062;
        finv_table[998] = 36'h034AB1068;
        finv_table[997] = 36'h036B8906C;
        finv_table[996] = 36'h038C6B071;
        finv_table[995] = 36'h03AD53073;
        finv_table[994] = 36'h03CE45078;
        finv_table[993] = 36'h03EF3F07C;
        finv_table[992] = 36'h041041081;
        finv_table[991] = 36'h04314B085;
        finv_table[990] = 36'h04525D088;
        finv_table[989] = 36'h04737908D;
        finv_table[988] = 36'h04949B090;
        finv_table[987] = 36'h04B5C7096;
        finv_table[986] = 36'h04D6FD09A;
        finv_table[985] = 36'h04F83909D;
        finv_table[984] = 36'h05197F0A2;
        finv_table[983] = 36'h053ACD0A6;
        finv_table[982] = 36'h055C230AA;
        finv_table[981] = 36'h057D810AF;
        finv_table[980] = 36'h059EE90B4;
        finv_table[979] = 36'h05C0590B7;
        finv_table[978] = 36'h05E1D10BC;
        finv_table[977] = 36'h0603530C0;
        finv_table[976] = 36'h0624DD0C4;
        finv_table[975] = 36'h06466F0C9;
        finv_table[974] = 36'h0668090CC;
        finv_table[973] = 36'h0689AD0D1;
        finv_table[972] = 36'h06AB590D5;
        finv_table[971] = 36'h06CD0D0DA;
        finv_table[970] = 36'h06EECB0DF;
        finv_table[969] = 36'h0710910E2;
        finv_table[968] = 36'h07325F0E7;
        finv_table[967] = 36'h0754370EC;
        finv_table[966] = 36'h0776170F0;
        finv_table[965] = 36'h0798010F4;
        finv_table[964] = 36'h07B9F10F9;
        finv_table[963] = 36'h07DBEB0FD;
        finv_table[962] = 36'h07FDEF102;
        finv_table[961] = 36'h081FFB105;
        finv_table[960] = 36'h08420F10A;
        finv_table[959] = 36'h08642D10F;
        finv_table[958] = 36'h088653112;
        finv_table[957] = 36'h08A883117;
        finv_table[956] = 36'h08CABB11C;
        finv_table[955] = 36'h08ECFB11F;
        finv_table[954] = 36'h090F45124;
        finv_table[953] = 36'h093197128;
        finv_table[952] = 36'h0953F312D;
        finv_table[951] = 36'h097657131;
        finv_table[950] = 36'h0998C5136;
        finv_table[949] = 36'h09BB3B13B;
        finv_table[948] = 36'h09DDB913E;
        finv_table[947] = 36'h0A0041144;
        finv_table[946] = 36'h0A22D3148;
        finv_table[945] = 36'h0A456D14C;
        finv_table[944] = 36'h0A680F150;
        finv_table[943] = 36'h0A8ABB156;
        finv_table[942] = 36'h0AAD7115B;
        finv_table[941] = 36'h0AD02F15E;
        finv_table[940] = 36'h0AF2F7163;
        finv_table[939] = 36'h0B15C7168;
        finv_table[938] = 36'h0B389F16B;
        finv_table[937] = 36'h0B5B83171;
        finv_table[936] = 36'h0B7E6D174;
        finv_table[935] = 36'h0BA16317A;
        finv_table[934] = 36'h0BC46117E;
        finv_table[933] = 36'h0BE767182;
        finv_table[932] = 36'h0C0A77188;
        finv_table[931] = 36'h0C2D9118C;
        finv_table[930] = 36'h0C50B3190;
        finv_table[929] = 36'h0C73DF195;
        finv_table[928] = 36'h0C971319A;
        finv_table[927] = 36'h0CBA5319F;
        finv_table[926] = 36'h0CDD991A2;
        finv_table[925] = 36'h0D00EB1A8;
        finv_table[924] = 36'h0D24451AC;
        finv_table[923] = 36'h0D47A71B0;
        finv_table[922] = 36'h0D6B151B6;
        finv_table[921] = 36'h0D8E8B1BB;
        finv_table[920] = 36'h0DB2091BE;
        finv_table[919] = 36'h0DD5931C4;
        finv_table[918] = 36'h0DF9251C9;
        finv_table[917] = 36'h0E1CBF1CC;
        finv_table[916] = 36'h0E40651D2;
        finv_table[915] = 36'h0E64131D6;
        finv_table[914] = 36'h0E87CB1DB;
        finv_table[913] = 36'h0EAB8B1DF;
        finv_table[912] = 36'h0ECF551E5;
        finv_table[911] = 36'h0EF3291EA;
        finv_table[910] = 36'h0F17071EF;
        finv_table[909] = 36'h0F3AEF1F3;
        finv_table[908] = 36'h0F5EDF1F8;
        finv_table[907] = 36'h0F82D91FC;
        finv_table[906] = 36'h0FA6DD201;
        finv_table[905] = 36'h0FCAE9205;
        finv_table[904] = 36'h0FEF0120B;
        finv_table[903] = 36'h101321210;
        finv_table[902] = 36'h10374B215;
        finv_table[901] = 36'h105B7D218;
        finv_table[900] = 36'h107FBB21F;
        finv_table[899] = 36'h10A401223;
        finv_table[898] = 36'h10C853228;
        finv_table[897] = 36'h10ECAD22D;
        finv_table[896] = 36'h111111232;
        finv_table[895] = 36'h11357D236;
        finv_table[894] = 36'h1159F523B;
        finv_table[893] = 36'h117E75240;
        finv_table[892] = 36'h11A301245;
        finv_table[891] = 36'h11C795249;
        finv_table[890] = 36'h11EC3324F;
        finv_table[889] = 36'h1210DB254;
        finv_table[888] = 36'h12358D259;
        finv_table[887] = 36'h125A4925E;
        finv_table[886] = 36'h127F0F262;
        finv_table[885] = 36'h12A3DF267;
        finv_table[884] = 36'h12C8B726B;
        finv_table[883] = 36'h12ED9B271;
        finv_table[882] = 36'h131287276;
        finv_table[881] = 36'h13377F27C;
        finv_table[880] = 36'h135C81280;
        finv_table[879] = 36'h13818B285;
        finv_table[878] = 36'h13A69F28A;
        finv_table[877] = 36'h13CBBF290;
        finv_table[876] = 36'h13F0E7294;
        finv_table[875] = 36'h14161B299;
        finv_table[874] = 36'h143B5729D;
        finv_table[873] = 36'h14609F2A3;
        finv_table[872] = 36'h1485EF2A8;
        finv_table[871] = 36'h14AB4B2AE;
        finv_table[870] = 36'h14D0B12B2;
        finv_table[869] = 36'h14F61F2B6;
        finv_table[868] = 36'h151B992BD;
        finv_table[867] = 36'h15411D2C1;
        finv_table[866] = 36'h1566AB2C6;
        finv_table[865] = 36'h158C432CB;
        finv_table[864] = 36'h15B1E52D0;
        finv_table[863] = 36'h15D7912D5;
        finv_table[862] = 36'h15FD492DB;
        finv_table[861] = 36'h1623092E1;
        finv_table[860] = 36'h1648D52E5;
        finv_table[859] = 36'h166EA92EB;
        finv_table[858] = 36'h1694892F0;
        finv_table[857] = 36'h16BA732F4;
        finv_table[856] = 36'h16E0672FA;
        finv_table[855] = 36'h1706672FF;
        finv_table[854] = 36'h172C6F303;
        finv_table[853] = 36'h175283309;
        finv_table[852] = 36'h1778A130E;
        finv_table[851] = 36'h179EC9313;
        finv_table[850] = 36'h17C4FB318;
        finv_table[849] = 36'h17EB3931E;
        finv_table[848] = 36'h181181324;
        finv_table[847] = 36'h1837D3329;
        finv_table[846] = 36'h185E2F32E;
        finv_table[845] = 36'h188495333;
        finv_table[844] = 36'h18AB07339;
        finv_table[843] = 36'h18D18333D;
        finv_table[842] = 36'h18F809343;
        finv_table[841] = 36'h191E9B349;
        finv_table[840] = 36'h19453734D;
        finv_table[839] = 36'h196BDD352;
        finv_table[838] = 36'h19928F358;
        finv_table[837] = 36'h19B94B35E;
        finv_table[836] = 36'h19E011363;
        finv_table[835] = 36'h1A06E1367;
        finv_table[834] = 36'h1A2DBD36E;
        finv_table[833] = 36'h1A54A3373;
        finv_table[832] = 36'h1A7B95379;
        finv_table[831] = 36'h1AA29137D;
        finv_table[830] = 36'h1AC997383;
        finv_table[829] = 36'h1AF0A9389;
        finv_table[828] = 36'h1B17C538E;
        finv_table[827] = 36'h1B3EED393;
        finv_table[826] = 36'h1B661F398;
        finv_table[825] = 36'h1B8D5B39D;
        finv_table[824] = 36'h1BB4A33A3;
        finv_table[823] = 36'h1BDBF53A8;
        finv_table[822] = 36'h1C03533AE;
        finv_table[821] = 36'h1C2ABB3B3;
        finv_table[820] = 36'h1C522F3B9;
        finv_table[819] = 36'h1C79AD3BE;
        finv_table[818] = 36'h1CA1373C4;
        finv_table[817] = 36'h1CC8CB3CA;
        finv_table[816] = 36'h1CF0693CE;
        finv_table[815] = 36'h1D18153D5;
        finv_table[814] = 36'h1D3FC93DA;
        finv_table[813] = 36'h1D67893E0;
        finv_table[812] = 36'h1D8F553E6;
        finv_table[811] = 36'h1DB72D3EB;
        finv_table[810] = 36'h1DDF0D3F0;
        finv_table[809] = 36'h1E06FB3F6;
        finv_table[808] = 36'h1E2EF33FB;
        finv_table[807] = 36'h1E56F5400;
        finv_table[806] = 36'h1E7F05407;
        finv_table[805] = 36'h1EA71D40B;
        finv_table[804] = 36'h1ECF43412;
        finv_table[803] = 36'h1EF773417;
        finv_table[802] = 36'h1F1FAF41D;
        finv_table[801] = 36'h1F47F5423;
        finv_table[800] = 36'h1F7047428;
        finv_table[799] = 36'h1F98A542E;
        finv_table[798] = 36'h1FC10D434;
        finv_table[797] = 36'h1FE981439;
        finv_table[796] = 36'h201201440;
        finv_table[795] = 36'h203A8B445;
        finv_table[794] = 36'h20632144A;
        finv_table[793] = 36'h208BC3450;
        finv_table[792] = 36'h20B46F455;
        finv_table[791] = 36'h20DD2945C;
        finv_table[790] = 36'h2105ED462;
        finv_table[789] = 36'h212EBB466;
        finv_table[788] = 36'h21579746D;
        finv_table[787] = 36'h21807D472;
        finv_table[786] = 36'h21A96F479;
        finv_table[785] = 36'h21D26D47F;
        finv_table[784] = 36'h21FB77484;
        finv_table[783] = 36'h22248D48A;
        finv_table[782] = 36'h224DAD490;
        finv_table[781] = 36'h2276D9495;
        finv_table[780] = 36'h22A01149B;
        finv_table[779] = 36'h22C9554A1;
        finv_table[778] = 36'h22F2A54A7;
        finv_table[777] = 36'h231BFF4AC;
        finv_table[776] = 36'h2345674B3;
        finv_table[775] = 36'h236ED94B8;
        finv_table[774] = 36'h2398574BF;
        finv_table[773] = 36'h23C1E34C5;
        finv_table[772] = 36'h23EB794CB;
        finv_table[771] = 36'h24151B4D1;
        finv_table[770] = 36'h243EC94D7;
        finv_table[769] = 36'h2468834DD;
        finv_table[768] = 36'h2492494E3;
        finv_table[767] = 36'h24BC194E8;
        finv_table[766] = 36'h24E5F74EF;
        finv_table[765] = 36'h250FE14F4;
        finv_table[764] = 36'h2539D74FA;
        finv_table[763] = 36'h2563D9500;
        finv_table[762] = 36'h258DE7507;
        finv_table[761] = 36'h25B80150D;
        finv_table[760] = 36'h25E227513;
        finv_table[759] = 36'h260C59519;
        finv_table[758] = 36'h26369751F;
        finv_table[757] = 36'h2660E1525;
        finv_table[756] = 36'h268B3752B;
        finv_table[755] = 36'h26B599530;
        finv_table[754] = 36'h26E009537;
        finv_table[753] = 36'h270A8353D;
        finv_table[752] = 36'h27350B543;
        finv_table[751] = 36'h275F9F54A;
        finv_table[750] = 36'h278A3D54F;
        finv_table[749] = 36'h27B4EB556;
        finv_table[748] = 36'h27DFA355C;
        finv_table[747] = 36'h280A67561;
        finv_table[746] = 36'h283539568;
        finv_table[745] = 36'h28601756F;
        finv_table[744] = 36'h288B01575;
        finv_table[743] = 36'h28B5F757B;
        finv_table[742] = 36'h28E0F9580;
        finv_table[741] = 36'h290C09587;
        finv_table[740] = 36'h29372558D;
        finv_table[739] = 36'h29624D593;
        finv_table[738] = 36'h298D8359B;
        finv_table[737] = 36'h29B8C35A1;
        finv_table[736] = 36'h29E4115A7;
        finv_table[735] = 36'h2A0F6D5AD;
        finv_table[734] = 36'h2A3AD35B3;
        finv_table[733] = 36'h2A66475BA;
        finv_table[732] = 36'h2A91C95C0;
        finv_table[731] = 36'h2ABD555C6;
        finv_table[730] = 36'h2AE8EF5CC;
        finv_table[729] = 36'h2B14975D3;
        finv_table[728] = 36'h2B40495D9;
        finv_table[727] = 36'h2B6C0B5E0;
        finv_table[726] = 36'h2B97D75E7;
        finv_table[725] = 36'h2BC3B15EC;
        finv_table[724] = 36'h2BEF975F2;
        finv_table[723] = 36'h2C1B8B5FA;
        finv_table[722] = 36'h2C478D600;
        finv_table[721] = 36'h2C7399607;
        finv_table[720] = 36'h2C9FB360D;
        finv_table[719] = 36'h2CCBDB613;
        finv_table[718] = 36'h2CF80F619;
        finv_table[717] = 36'h2D2451620;
        finv_table[716] = 36'h2D509F626;
        finv_table[715] = 36'h2D7CFB62D;
        finv_table[714] = 36'h2DA963634;
        finv_table[713] = 36'h2DD5D963B;
        finv_table[712] = 36'h2E025B641;
        finv_table[711] = 36'h2E2EEB647;
        finv_table[710] = 36'h2E5B8764D;
        finv_table[709] = 36'h2E8831655;
        finv_table[708] = 36'h2EB4E965B;
        finv_table[707] = 36'h2EE1AD661;
        finv_table[706] = 36'h2F0E7F668;
        finv_table[705] = 36'h2F3B5F66F;
        finv_table[704] = 36'h2F684B676;
        finv_table[703] = 36'h2F954567D;
        finv_table[702] = 36'h2FC24B682;
        finv_table[701] = 36'h2FEF5F68A;
        finv_table[700] = 36'h301C81691;
        finv_table[699] = 36'h3049B1697;
        finv_table[698] = 36'h3076ED69D;
        finv_table[697] = 36'h30A4376A4;
        finv_table[696] = 36'h30D18F6AB;
        finv_table[695] = 36'h30FEF56B3;
        finv_table[694] = 36'h312C676B9;
        finv_table[693] = 36'h3159E76C0;
        finv_table[692] = 36'h3187756C7;
        finv_table[691] = 36'h31B50F6CC;
        finv_table[690] = 36'h31E2B96D4;
        finv_table[689] = 36'h32106F6DA;
        finv_table[688] = 36'h323E336E1;
        finv_table[687] = 36'h326C056E8;
        finv_table[686] = 36'h3299E56EF;
        finv_table[685] = 36'h32C7D36F6;
        finv_table[684] = 36'h32F5CD6FC;
        finv_table[683] = 36'h3323D7704;
        finv_table[682] = 36'h3351ED70A;
        finv_table[681] = 36'h338013712;
        finv_table[680] = 36'h33AE45719;
        finv_table[679] = 36'h33DC85720;
        finv_table[678] = 36'h340AD3726;
        finv_table[677] = 36'h34392F72D;
        finv_table[676] = 36'h346799734;
        finv_table[675] = 36'h34961173C;
        finv_table[674] = 36'h34C499743;
        finv_table[673] = 36'h34F32D74A;
        finv_table[672] = 36'h3521CF751;
        finv_table[671] = 36'h35507F758;
        finv_table[670] = 36'h357F3D75E;
        finv_table[669] = 36'h35AE0B766;
        finv_table[668] = 36'h35DCE576D;
        finv_table[667] = 36'h360BCD773;
        finv_table[666] = 36'h363AC577B;
        finv_table[665] = 36'h3669CB783;
        finv_table[664] = 36'h3698DF78A;
        finv_table[663] = 36'h36C801791;
        finv_table[662] = 36'h36F731798;
        finv_table[661] = 36'h37266F79F;
        finv_table[660] = 36'h3755BD7A7;
        finv_table[659] = 36'h3785177AD;
        finv_table[658] = 36'h37B4817B4;
        finv_table[657] = 36'h37E3F97BB;
        finv_table[656] = 36'h3813817C3;
        finv_table[655] = 36'h3843157CA;
        finv_table[654] = 36'h3872B97D1;
        finv_table[653] = 36'h38A26B7D8;
        finv_table[652] = 36'h38D22D7E1;
        finv_table[651] = 36'h3901FB7E7;
        finv_table[650] = 36'h3931D97EE;
        finv_table[649] = 36'h3961C77F6;
        finv_table[648] = 36'h3991C17FD;
        finv_table[647] = 36'h39C1CB804;
        finv_table[646] = 36'h39F1E580C;
        finv_table[645] = 36'h3A220D814;
        finv_table[644] = 36'h3A524381B;
        finv_table[643] = 36'h3A8287822;
        finv_table[642] = 36'h3AB2DB829;
        finv_table[641] = 36'h3AE33F831;
        finv_table[640] = 36'h3B13B1839;
        finv_table[639] = 36'h3B4431840;
        finv_table[638] = 36'h3B74C1848;
        finv_table[637] = 36'h3BA55F84F;
        finv_table[636] = 36'h3BD60D857;
        finv_table[635] = 36'h3C06C985E;
        finv_table[634] = 36'h3C3795866;
        finv_table[633] = 36'h3C686F86C;
        finv_table[632] = 36'h3C9959874;
        finv_table[631] = 36'h3CCA5387D;
        finv_table[630] = 36'h3CFB5B884;
        finv_table[629] = 36'h3D2C7188B;
        finv_table[628] = 36'h3D5D99894;
        finv_table[627] = 36'h3D8ECD89A;
        finv_table[626] = 36'h3DC0138A2;
        finv_table[625] = 36'h3DF1678AA;
        finv_table[624] = 36'h3E22CB8B2;
        finv_table[623] = 36'h3E543D8B8;
        finv_table[622] = 36'h3E85C18C1;
        finv_table[621] = 36'h3EB7518C8;
        finv_table[620] = 36'h3EE8F38D0;
        finv_table[619] = 36'h3F1AA38D7;
        finv_table[618] = 36'h3F4C658E0;
        finv_table[617] = 36'h3F7E338E7;
        finv_table[616] = 36'h3FB0138EF;
        finv_table[615] = 36'h3FE2018F6;
        finv_table[614] = 36'h4014018FF;
        finv_table[613] = 36'h40460F907;
        finv_table[612] = 36'h40782D90F;
        finv_table[611] = 36'h40AA59916;
        finv_table[610] = 36'h40DC9791E;
        finv_table[609] = 36'h410EE3926;
        finv_table[608] = 36'h41414192F;
        finv_table[607] = 36'h4173AD936;
        finv_table[606] = 36'h41A62993E;
        finv_table[605] = 36'h41D8B5945;
        finv_table[604] = 36'h420B5194D;
        finv_table[603] = 36'h423DFD955;
        finv_table[602] = 36'h4270B995D;
        finv_table[601] = 36'h42A385965;
        finv_table[600] = 36'h42D66196D;
        finv_table[599] = 36'h43094D975;
        finv_table[598] = 36'h433C4997D;
        finv_table[597] = 36'h436F55985;
        finv_table[596] = 36'h43A27398F;
        finv_table[595] = 36'h43D59F996;
        finv_table[594] = 36'h4408DB99E;
        finv_table[593] = 36'h443C299A7;
        finv_table[592] = 36'h446F859AE;
        finv_table[591] = 36'h44A2F39B7;
        finv_table[590] = 36'h44D6719BF;
        finv_table[589] = 36'h4509FF9C7;
        finv_table[588] = 36'h453D9D9CF;
        finv_table[587] = 36'h45714D9D8;
        finv_table[586] = 36'h45A50B9DF;
        finv_table[585] = 36'h45D8DB9E7;
        finv_table[584] = 36'h460CBB9EF;
        finv_table[583] = 36'h4640AD9F9;
        finv_table[582] = 36'h4674ADA00;
        finv_table[581] = 36'h46A8BFA08;
        finv_table[580] = 36'h46DCE3A12;
        finv_table[579] = 36'h471115A19;
        finv_table[578] = 36'h474559A21;
        finv_table[577] = 36'h4779AFA2B;
        finv_table[576] = 36'h47AE13A32;
        finv_table[575] = 36'h47E289A3A;
        finv_table[574] = 36'h481711A43;
        finv_table[573] = 36'h484BA9A4C;
        finv_table[572] = 36'h488051A54;
        finv_table[571] = 36'h48B50BA5D;
        finv_table[570] = 36'h48E9D5A65;
        finv_table[569] = 36'h491EB1A6E;
        finv_table[568] = 36'h49539DA76;
        finv_table[567] = 36'h49889BA7F;
        finv_table[566] = 36'h49BDA9A87;
        finv_table[565] = 36'h49F2C9A90;
        finv_table[564] = 36'h4A27F9A97;
        finv_table[563] = 36'h4A5D3BAA0;
        finv_table[562] = 36'h4A928FAA9;
        finv_table[561] = 36'h4AC7F3AB2;
        finv_table[560] = 36'h4AFD69ABB;
        finv_table[559] = 36'h4B32EFAC2;
        finv_table[558] = 36'h4B6889ACD;
        finv_table[557] = 36'h4B9E31AD4;
        finv_table[556] = 36'h4BD3EDADD;
        finv_table[555] = 36'h4C09B9AE6;
        finv_table[554] = 36'h4C3F97AEF;
        finv_table[553] = 36'h4C7587AF8;
        finv_table[552] = 36'h4CAB87B00;
        finv_table[551] = 36'h4CE199B08;
        finv_table[550] = 36'h4D17BDB11;
        finv_table[549] = 36'h4D4DF3B1A;
        finv_table[548] = 36'h4D843BB23;
        finv_table[547] = 36'h4DBA93B2C;
        finv_table[546] = 36'h4DF0FFB35;
        finv_table[545] = 36'h4E277BB3E;
        finv_table[544] = 36'h4E5E09B47;
        finv_table[543] = 36'h4E94A9B4F;
        finv_table[542] = 36'h4ECB5BB58;
        finv_table[541] = 36'h4F021FB61;
        finv_table[540] = 36'h4F38F5B6B;
        finv_table[539] = 36'h4F6FDDB74;
        finv_table[538] = 36'h4FA6D7B7D;
        finv_table[537] = 36'h4FDDE3B86;
        finv_table[536] = 36'h501501B8F;
        finv_table[535] = 36'h504C31B98;
        finv_table[534] = 36'h508373BA1;
        finv_table[533] = 36'h50BAC7BAA;
        finv_table[532] = 36'h50F22DBB3;
        finv_table[531] = 36'h5129A5BBC;
        finv_table[530] = 36'h516131BC6;
        finv_table[529] = 36'h5198CFBCF;
        finv_table[528] = 36'h51D07DBD7;
        finv_table[527] = 36'h52083FBE0;
        finv_table[526] = 36'h524015BEB;
        finv_table[525] = 36'h5277FBBF3;
        finv_table[524] = 36'h52AFF5BFD;
        finv_table[523] = 36'h52E801C06;
        finv_table[522] = 36'h53201FC0F;
        finv_table[521] = 36'h53584FC18;
        finv_table[520] = 36'h539093C21;
        finv_table[519] = 36'h53C8E9C2A;
        finv_table[518] = 36'h540153C34;
        finv_table[517] = 36'h5439CFC3E;
        finv_table[516] = 36'h54725DC47;
        finv_table[515] = 36'h54AAFFC51;
        finv_table[514] = 36'h54E3B3C5A;
        finv_table[513] = 36'h551C7BC64;
        finv_table[512] = 36'h555553C6C;
        finv_table[511] = 36'h558E41C76;
        finv_table[510] = 36'h55C741C80;
        finv_table[509] = 36'h560055C8A;
        finv_table[508] = 36'h56397BC93;
        finv_table[507] = 36'h5672B3C9C;
        finv_table[506] = 36'h56AC01CA7;
        finv_table[505] = 36'h56E55FCAF;
        finv_table[504] = 36'h571ED3CBA;
        finv_table[503] = 36'h575859CC3;
        finv_table[502] = 36'h5791F3CCD;
        finv_table[501] = 36'h57CB9FCD6;
        finv_table[500] = 36'h58055FCE0;
        finv_table[499] = 36'h583F33CEA;
        finv_table[498] = 36'h587919CF3;
        finv_table[497] = 36'h58B315CFE;
        finv_table[496] = 36'h58ED23D08;
        finv_table[495] = 36'h592743D10;
        finv_table[494] = 36'h596179D1B;
        finv_table[493] = 36'h599BC1D24;
        finv_table[492] = 36'h59D61FD2F;
        finv_table[491] = 36'h5A108FD39;
        finv_table[490] = 36'h5A4B11D41;
        finv_table[489] = 36'h5A85A9D4B;
        finv_table[488] = 36'h5AC055D55;
        finv_table[487] = 36'h5AFB15D60;
        finv_table[486] = 36'h5B35E9D6A;
        finv_table[485] = 36'h5B70CFD73;
        finv_table[484] = 36'h5BABCBD7D;
        finv_table[483] = 36'h5BE6DBD88;
        finv_table[482] = 36'h5C21FFD92;
        finv_table[481] = 36'h5C5D35D9B;
        finv_table[480] = 36'h5C9881DA5;
        finv_table[479] = 36'h5CD3E1DAF;
        finv_table[478] = 36'h5D0F55DB9;
        finv_table[477] = 36'h5D4ADFDC5;
        finv_table[476] = 36'h5D867BDCE;
        finv_table[475] = 36'h5DC22DDD9;
        finv_table[474] = 36'h5DFDF1DE2;
        finv_table[473] = 36'h5E39CDDEE;
        finv_table[472] = 36'h5E75BBDF8;
        finv_table[471] = 36'h5EB1BDE01;
        finv_table[470] = 36'h5EEDD5E0C;
        finv_table[469] = 36'h5F2A01E16;
        finv_table[468] = 36'h5F6643E21;
        finv_table[467] = 36'h5FA297E2A;
        finv_table[466] = 36'h5FDF03E36;
        finv_table[465] = 36'h601B7FE3E;
        finv_table[464] = 36'h605815E4A;
        finv_table[463] = 36'h6094BDE54;
        finv_table[462] = 36'h60D17BE5F;
        finv_table[461] = 36'h610E4DE69;
        finv_table[460] = 36'h614B35E73;
        finv_table[459] = 36'h618833E7F;
        finv_table[458] = 36'h61C543E88;
        finv_table[457] = 36'h62026BE94;
        finv_table[456] = 36'h623FA5E9D;
        finv_table[455] = 36'h627CF7EA8;
        finv_table[454] = 36'h62BA5DEB3;
        finv_table[453] = 36'h62F7D9EBD;
        finv_table[452] = 36'h63356BEC9;
        finv_table[451] = 36'h637311ED3;
        finv_table[450] = 36'h63B0CDEDE;
        finv_table[449] = 36'h63EE9DEE8;
        finv_table[448] = 36'h642C85EF4;
        finv_table[447] = 36'h646A81EFE;
        finv_table[446] = 36'h64A893F09;
        finv_table[445] = 36'h64E6B9F13;
        finv_table[444] = 36'h6524F7F1E;
        finv_table[443] = 36'h65634BF2A;
        finv_table[442] = 36'h65A1B1F33;
        finv_table[441] = 36'h65E031F3F;
        finv_table[440] = 36'h661EC5F4A;
        finv_table[439] = 36'h665D6FF55;
        finv_table[438] = 36'h669C31F61;
        finv_table[437] = 36'h66DB07F6C;
        finv_table[436] = 36'h6719F1F75;
        finv_table[435] = 36'h6758F3F80;
        finv_table[434] = 36'h67980DF8C;
        finv_table[433] = 36'h67D73BF97;
        finv_table[432] = 36'h681681FA3;
        finv_table[431] = 36'h6855DBFAD;
        finv_table[430] = 36'h68954DFB9;
        finv_table[429] = 36'h68D4D3FC3;
        finv_table[428] = 36'h691471FCE;
        finv_table[427] = 36'h695427FDA;
        finv_table[426] = 36'h6993F1FE5;
        finv_table[425] = 36'h69D3D3FF0;
        finv_table[424] = 36'h6A13CDFFD;
        finv_table[423] = 36'h6A53DB004;
        finv_table[422] = 36'h6A93FF009;
        finv_table[421] = 36'h6AD43B00F;
        finv_table[420] = 36'h6B148D014;
        finv_table[419] = 36'h6B54F701A;
        finv_table[418] = 36'h6B9579020;
        finv_table[417] = 36'h6BD60F025;
        finv_table[416] = 36'h6C16C102C;
        finv_table[415] = 36'h6C5785031;
        finv_table[414] = 36'h6C9861037;
        finv_table[413] = 36'h6CD95503D;
        finv_table[412] = 36'h6D1A5F042;
        finv_table[411] = 36'h6D5B81048;
        finv_table[410] = 36'h6D9CBB04E;
        finv_table[409] = 36'h6DDE0D054;
        finv_table[408] = 36'h6E1F7505A;
        finv_table[407] = 36'h6E60F5060;
        finv_table[406] = 36'h6EA28B066;
        finv_table[405] = 36'h6EE43B06C;
        finv_table[404] = 36'h6F25FF071;
        finv_table[403] = 36'h6F67DD077;
        finv_table[402] = 36'h6FA9D107D;
        finv_table[401] = 36'h6FEBDF083;
        finv_table[400] = 36'h702E03089;
        finv_table[399] = 36'h70704108F;
        finv_table[398] = 36'h70B295095;
        finv_table[397] = 36'h70F50109B;
        finv_table[396] = 36'h7137850A1;
        finv_table[395] = 36'h717A210A7;
        finv_table[394] = 36'h71BCD50AD;
        finv_table[393] = 36'h71FFA10B3;
        finv_table[392] = 36'h7242850B9;
        finv_table[391] = 36'h7285830BF;
        finv_table[390] = 36'h72C8970C5;
        finv_table[389] = 36'h730BC50CB;
        finv_table[388] = 36'h734F090D1;
        finv_table[387] = 36'h7392670D7;
        finv_table[386] = 36'h73D5DD0DD;
        finv_table[385] = 36'h74196F0E4;
        finv_table[384] = 36'h745D150EA;
        finv_table[383] = 36'h74A0D50F0;
        finv_table[382] = 36'h74E4AD0F6;
        finv_table[381] = 36'h75289F0FC;
        finv_table[380] = 36'h756CA9102;
        finv_table[379] = 36'h75B0CD109;
        finv_table[378] = 36'h75F50910F;
        finv_table[377] = 36'h76395D115;
        finv_table[376] = 36'h767DCB11B;
        finv_table[375] = 36'h76C253122;
        finv_table[374] = 36'h7706F3128;
        finv_table[373] = 36'h774BAB12E;
        finv_table[372] = 36'h77907F135;
        finv_table[371] = 36'h77D56913A;
        finv_table[370] = 36'h781A6F141;
        finv_table[369] = 36'h785F8D147;
        finv_table[368] = 36'h78A4C714E;
        finv_table[367] = 36'h78EA17154;
        finv_table[366] = 36'h792F8115A;
        finv_table[365] = 36'h797507161;
        finv_table[364] = 36'h79BAA3167;
        finv_table[363] = 36'h7A005D16E;
        finv_table[362] = 36'h7A462D174;
        finv_table[361] = 36'h7A8C1917B;
        finv_table[360] = 36'h7AD21D181;
        finv_table[359] = 36'h7B183D188;
        finv_table[358] = 36'h7B5E7518E;
        finv_table[357] = 36'h7BA4CB195;
        finv_table[356] = 36'h7BEB3719B;
        finv_table[355] = 36'h7C31BD1A1;
        finv_table[354] = 36'h7C785F1A8;
        finv_table[353] = 36'h7CBF1B1AF;
        finv_table[352] = 36'h7D05F11B5;
        finv_table[351] = 36'h7D4CE31BC;
        finv_table[350] = 36'h7D93ED1C3;
        finv_table[349] = 36'h7DDB131C9;
        finv_table[348] = 36'h7E22531D0;
        finv_table[347] = 36'h7E69AF1D7;
        finv_table[346] = 36'h7EB1211DD;
        finv_table[345] = 36'h7EF8B31E4;
        finv_table[344] = 36'h7F405F1EB;
        finv_table[343] = 36'h7F88231F1;
        finv_table[342] = 36'h7FD0031F8;
        finv_table[341] = 36'h8017FF1FF;
        finv_table[340] = 36'h806015205;
        finv_table[339] = 36'h80A84720C;
        finv_table[338] = 36'h80F093213;
        finv_table[337] = 36'h8138FB21A;
        finv_table[336] = 36'h81817F221;
        finv_table[335] = 36'h81CA1D227;
        finv_table[334] = 36'h8212D722E;
        finv_table[333] = 36'h825BAD235;
        finv_table[332] = 36'h82A49D23C;
        finv_table[331] = 36'h82EDA9243;
        finv_table[330] = 36'h8336D324A;
        finv_table[329] = 36'h838015251;
        finv_table[328] = 36'h83C975258;
        finv_table[327] = 36'h8412EF25E;
        finv_table[326] = 36'h845C89266;
        finv_table[325] = 36'h84A63B26D;
        finv_table[324] = 36'h84F00B274;
        finv_table[323] = 36'h8539F527B;
        finv_table[322] = 36'h8583FB281;
        finv_table[321] = 36'h85CE1F289;
        finv_table[320] = 36'h86185F290;
        finv_table[319] = 36'h8662BB297;
        finv_table[318] = 36'h86AD3329E;
        finv_table[317] = 36'h86F7C72A5;
        finv_table[316] = 36'h8742792AC;
        finv_table[315] = 36'h878D472B3;
        finv_table[314] = 36'h87D8312BA;
        finv_table[313] = 36'h8823392C2;
        finv_table[312] = 36'h886E5D2C9;
        finv_table[311] = 36'h88B99D2D0;
        finv_table[310] = 36'h8904FB2D7;
        finv_table[309] = 36'h8950752DE;
        finv_table[308] = 36'h899C0D2E6;
        finv_table[307] = 36'h89E7C12ED;
        finv_table[306] = 36'h8A33932F4;
        finv_table[305] = 36'h8A7F812FB;
        finv_table[304] = 36'h8ACB8F303;
        finv_table[303] = 36'h8B17B730A;
        finv_table[302] = 36'h8B63FF312;
        finv_table[301] = 36'h8BB063319;
        finv_table[300] = 36'h8BFCE5320;
        finv_table[299] = 36'h8C4985328;
        finv_table[298] = 36'h8C964132F;
        finv_table[297] = 36'h8CE31D337;
        finv_table[296] = 36'h8D301533E;
        finv_table[295] = 36'h8D7D2D346;
        finv_table[294] = 36'h8DCA6134D;
        finv_table[293] = 36'h8E17B3354;
        finv_table[292] = 36'h8E652535C;
        finv_table[291] = 36'h8EB2B3363;
        finv_table[290] = 36'h8F006136B;
        finv_table[289] = 36'h8F4E2D373;
        finv_table[288] = 36'h8F9C1537A;
        finv_table[287] = 36'h8FEA1F382;
        finv_table[286] = 36'h903845389;
        finv_table[285] = 36'h90868B391;
        finv_table[284] = 36'h90D4EF399;
        finv_table[283] = 36'h9123713A0;
        finv_table[282] = 36'h9172133A8;
        finv_table[281] = 36'h91C0D33B0;
        finv_table[280] = 36'h920FB33B8;
        finv_table[279] = 36'h925EAF3BF;
        finv_table[278] = 36'h92ADCD3C7;
        finv_table[277] = 36'h92FD093CF;
        finv_table[276] = 36'h934C653D7;
        finv_table[275] = 36'h939BDF3DE;
        finv_table[274] = 36'h93EB7B3E7;
        finv_table[273] = 36'h943B333EE;
        finv_table[272] = 36'h948B0D3F6;
        finv_table[271] = 36'h94DB053FE;
        finv_table[270] = 36'h952B1D406;
        finv_table[269] = 36'h957B5540E;
        finv_table[268] = 36'h95CBAD416;
        finv_table[267] = 36'h961C2541E;
        finv_table[266] = 36'h966CBD426;
        finv_table[265] = 36'h96BD7542E;
        finv_table[264] = 36'h970E4D436;
        finv_table[263] = 36'h975F4543E;
        finv_table[262] = 36'h97B05D446;
        finv_table[261] = 36'h98019544E;
        finv_table[260] = 36'h9852ED456;
        finv_table[259] = 36'h98A46745E;
        finv_table[258] = 36'h98F601466;
        finv_table[257] = 36'h9947BB46E;
        finv_table[256] = 36'h999997477;
        finv_table[255] = 36'h99EB9347F;
        finv_table[254] = 36'h9A3DAF487;
        finv_table[253] = 36'h9A8FED48F;
        finv_table[252] = 36'h9AE24B497;
        finv_table[251] = 36'h9B34CB4A0;
        finv_table[250] = 36'h9B876D4A8;
        finv_table[249] = 36'h9BDA2F4B0;
        finv_table[248] = 36'h9C2D134B9;
        finv_table[247] = 36'h9C80174C1;
        finv_table[246] = 36'h9CD33D4C9;
        finv_table[245] = 36'h9D26854D2;
        finv_table[244] = 36'h9D79EF4DA;
        finv_table[243] = 36'h9DCD794E2;
        finv_table[242] = 36'h9E21274EB;
        finv_table[241] = 36'h9E74F54F3;
        finv_table[240] = 36'h9EC8E74FC;
        finv_table[239] = 36'h9F1CF9504;
        finv_table[238] = 36'h9F712F50D;
        finv_table[237] = 36'h9FC585515;
        finv_table[236] = 36'hA019FF51E;
        finv_table[235] = 36'hA06E9B527;
        finv_table[234] = 36'hA0C35952F;
        finv_table[233] = 36'hA11839538;
        finv_table[232] = 36'hA16D3D541;
        finv_table[231] = 36'hA1C263549;
        finv_table[230] = 36'hA217AB552;
        finv_table[229] = 36'hA26D1755B;
        finv_table[228] = 36'hA2C2A5563;
        finv_table[227] = 36'hA3185756C;
        finv_table[226] = 36'hA36E2B575;
        finv_table[225] = 36'hA3C42357E;
        finv_table[224] = 36'hA41A3F587;
        finv_table[223] = 36'hA4707D58F;
        finv_table[222] = 36'hA4C6DF598;
        finv_table[221] = 36'hA51D655A1;
        finv_table[220] = 36'hA5740D5AA;
        finv_table[219] = 36'hA5CADB5B3;
        finv_table[218] = 36'hA621CB5BC;
        finv_table[217] = 36'hA678DF5C5;
        finv_table[216] = 36'hA6D0175CE;
        finv_table[215] = 36'hA727735D7;
        finv_table[214] = 36'hA77EF55E0;
        finv_table[213] = 36'hA7D6995E9;
        finv_table[212] = 36'hA82E635F2;
        finv_table[211] = 36'hA8864F5FB;
        finv_table[210] = 36'hA8DE61604;
        finv_table[209] = 36'hA9369960E;
        finv_table[208] = 36'hA98EF3617;
        finv_table[207] = 36'hA9E773620;
        finv_table[206] = 36'hAA4017629;
        finv_table[205] = 36'hAA98E1632;
        finv_table[204] = 36'hAAF1CF63B;
        finv_table[203] = 36'hAB4AE3645;
        finv_table[202] = 36'hABA41D64E;
        finv_table[201] = 36'hABFD7B657;
        finv_table[200] = 36'hAC56FF661;
        finv_table[199] = 36'hACB0A766A;
        finv_table[198] = 36'hAD0A77674;
        finv_table[197] = 36'hAD646B67D;
        finv_table[196] = 36'hADBE85686;
        finv_table[195] = 36'hAE18C5690;
        finv_table[194] = 36'hAE732B699;
        finv_table[193] = 36'hAECDB76A3;
        finv_table[192] = 36'hAF28696AC;
        finv_table[191] = 36'hAF83416B6;
        finv_table[190] = 36'hAFDE3F6BF;
        finv_table[189] = 36'hB039656C9;
        finv_table[188] = 36'hB094B16D3;
        finv_table[187] = 36'hB0F0236DD;
        finv_table[186] = 36'hB14BBB6E6;
        finv_table[185] = 36'hB1A77B6F0;
        finv_table[184] = 36'hB203616F9;
        finv_table[183] = 36'hB25F6F703;
        finv_table[182] = 36'hB2BBA370D;
        finv_table[181] = 36'hB317FF717;
        finv_table[180] = 36'hB37481720;
        finv_table[179] = 36'hB3D12D72B;
        finv_table[178] = 36'hB42DFD734;
        finv_table[177] = 36'hB48AF773E;
        finv_table[176] = 36'hB4E819748;
        finv_table[175] = 36'hB54561752;
        finv_table[174] = 36'hB5A2D175C;
        finv_table[173] = 36'hB6006B766;
        finv_table[172] = 36'hB65E2B770;
        finv_table[171] = 36'hB6BC1577A;
        finv_table[170] = 36'hB71A25784;
        finv_table[169] = 36'hB7785F78E;
        finv_table[168] = 36'hB7D6C1798;
        finv_table[167] = 36'hB8354B7A2;
        finv_table[166] = 36'hB893FF7AD;
        finv_table[165] = 36'hB8F2DB7B7;
        finv_table[164] = 36'hB951DF7C1;
        finv_table[163] = 36'hB9B10D7CB;
        finv_table[162] = 36'hBA10657D6;
        finv_table[161] = 36'hBA6FE57E0;
        finv_table[160] = 36'hBACF8F7EA;
        finv_table[159] = 36'hBB2F617F4;
        finv_table[158] = 36'hBB8F5D7FF;
        finv_table[157] = 36'hBBEF83809;
        finv_table[156] = 36'hBC4FD3814;
        finv_table[155] = 36'hBCB04D81E;
        finv_table[154] = 36'hBD10F1829;
        finv_table[153] = 36'hBD71BD833;
        finv_table[152] = 36'hBDD2B583E;
        finv_table[151] = 36'hBE33D7848;
        finv_table[150] = 36'hBE9523853;
        finv_table[149] = 36'hBEF69B85E;
        finv_table[148] = 36'hBF583B868;
        finv_table[147] = 36'hBFBA07873;
        finv_table[146] = 36'hC01BFF87E;
        finv_table[145] = 36'hC07E21888;
        finv_table[144] = 36'hC0E06D893;
        finv_table[143] = 36'hC142E589E;
        finv_table[142] = 36'hC1A5898A9;
        finv_table[141] = 36'hC208558B3;
        finv_table[140] = 36'hC26B518BE;
        finv_table[139] = 36'hC2CE758C9;
        finv_table[138] = 36'hC331C78D4;
        finv_table[137] = 36'hC395458DF;
        finv_table[136] = 36'hC3F8ED8EA;
        finv_table[135] = 36'hC45CC38F5;
        finv_table[134] = 36'hC4C0C3900;
        finv_table[133] = 36'hC524F190B;
        finv_table[132] = 36'hC58949916;
        finv_table[131] = 36'hC5EDCF921;
        finv_table[130] = 36'hC6528592D;
        finv_table[129] = 36'hC6B763938;
        finv_table[128] = 36'hC71C6F943;
        finv_table[127] = 36'hC781A794E;
        finv_table[126] = 36'hC7E70F95A;
        finv_table[125] = 36'hC84CA1964;
        finv_table[124] = 36'hC8B263970;
        finv_table[123] = 36'hC9185197B;
        finv_table[122] = 36'hC97E6D987;
        finv_table[121] = 36'hC9E4B5992;
        finv_table[120] = 36'hCA4B2D99E;
        finv_table[119] = 36'hCAB1D39A9;
        finv_table[118] = 36'hCB18A59B4;
        finv_table[117] = 36'hCB7FA79C0;
        finv_table[116] = 36'hCBE6D79CC;
        finv_table[115] = 36'hCC4E339D7;
        finv_table[114] = 36'hCCB5C19E3;
        finv_table[113] = 36'hCD1D7B9EE;
        finv_table[112] = 36'hCD85659FA;
        finv_table[111] = 36'hCDED7FA06;
        finv_table[110] = 36'hCE55C5A11;
        finv_table[109] = 36'hCEBE3DA1E;
        finv_table[108] = 36'hCF26E1A29;
        finv_table[107] = 36'hCF8FB7A35;
        finv_table[106] = 36'hCFF8BDA41;
        finv_table[105] = 36'hD061F1A4D;
        finv_table[104] = 36'hD0CB55A59;
        finv_table[103] = 36'hD134EBA65;
        finv_table[102] = 36'hD19EAFA71;
        finv_table[101] = 36'hD208A3A7D;
        finv_table[100] = 36'hD272C7A89;
        finv_table[99] = 36'hD2DD1BA95;
        finv_table[98] = 36'hD347A1AA1;
        finv_table[97] = 36'hD3B257AAD;
        finv_table[96] = 36'hD41D3FABA;
        finv_table[95] = 36'hD48857AC6;
        finv_table[94] = 36'hD4F39FAD2;
        finv_table[93] = 36'hD55F19ADE;
        finv_table[92] = 36'hD5CAC5AEB;
        finv_table[91] = 36'hD636A1AF7;
        finv_table[90] = 36'hD6A2B1B04;
        finv_table[89] = 36'hD70EF1B10;
        finv_table[88] = 36'hD77B61B1C;
        finv_table[87] = 36'hD7E807B29;
        finv_table[86] = 36'hD854DBB35;
        finv_table[85] = 36'hD8C1E5B42;
        finv_table[84] = 36'hD92F1DB4E;
        finv_table[83] = 36'hD99C8BB5B;
        finv_table[82] = 36'hDA0A2BB68;
        finv_table[81] = 36'hDA77FFB75;
        finv_table[80] = 36'hDAE603B81;
        finv_table[79] = 36'hDB543DB8E;
        finv_table[78] = 36'hDBC2A9B9B;
        finv_table[77] = 36'hDC3149BA8;
        finv_table[76] = 36'hDCA019BB4;
        finv_table[75] = 36'hDD0F1FBC1;
        finv_table[74] = 36'hDD7E59BCE;
        finv_table[73] = 36'hDDEDC7BDB;
        finv_table[72] = 36'hDE5D69BE8;
        finv_table[71] = 36'hDECD3FBF5;
        finv_table[70] = 36'hDF3D4DC03;
        finv_table[69] = 36'hDFAD8BC10;
        finv_table[68] = 36'hE01DFFC1D;
        finv_table[67] = 36'hE08EA7C2A;
        finv_table[66] = 36'hE0FF83C37;
        finv_table[65] = 36'hE17095C44;
        finv_table[64] = 36'hE1E1DFC52;
        finv_table[63] = 36'hE2535BC5F;
        finv_table[62] = 36'hE2C50FC6D;
        finv_table[61] = 36'hE336F5C7A;
        finv_table[60] = 36'hE3A913C87;
        finv_table[59] = 36'hE41B67C95;
        finv_table[58] = 36'hE48DF1CA2;
        finv_table[57] = 36'hE500B1CB0;
        finv_table[56] = 36'hE573A7CBD;
        finv_table[55] = 36'hE5E6D5CCB;
        finv_table[54] = 36'hE65A39CD9;
        finv_table[53] = 36'hE6CDD3CE6;
        finv_table[52] = 36'hE741A5CF4;
        finv_table[51] = 36'hE7B5AFD02;
        finv_table[50] = 36'hE829EFD10;
        finv_table[49] = 36'hE89E67D1E;
        finv_table[48] = 36'hE91315D2B;
        finv_table[47] = 36'hE987FFD3A;
        finv_table[46] = 36'hE9FD1DD48;
        finv_table[45] = 36'hEA7275D56;
        finv_table[44] = 36'hEAE803D64;
        finv_table[43] = 36'hEB5DCBD72;
        finv_table[42] = 36'hEBD3CBD80;
        finv_table[41] = 36'hEC4A05D8E;
        finv_table[40] = 36'hECC077D9C;
        finv_table[39] = 36'hED3721DAA;
        finv_table[38] = 36'hEDAE07DB9;
        finv_table[37] = 36'hEE2523DC7;
        finv_table[36] = 36'hEE9C7BDD6;
        finv_table[35] = 36'hEF140BDE4;
        finv_table[34] = 36'hEF8BD7DF3;
        finv_table[33] = 36'hF003DBE01;
        finv_table[32] = 36'hF07C1BE10;
        finv_table[31] = 36'hF0F493E1E;
        finv_table[30] = 36'hF16D49E2D;
        finv_table[29] = 36'hF1E635E3B;
        finv_table[28] = 36'hF25F5FE4A;
        finv_table[27] = 36'hF2D8C5E59;
        finv_table[26] = 36'hF35265E68;
        finv_table[25] = 36'hF3CC3FE77;
        finv_table[24] = 36'hF44655E85;
        finv_table[23] = 36'hF4C0A7E94;
        finv_table[22] = 36'hF53B35EA3;
        finv_table[21] = 36'hF5B5FFEB2;
        finv_table[20] = 36'hF63105EC1;
        finv_table[19] = 36'hF6AC49ED1;
        finv_table[18] = 36'hF727C7EDF;
        finv_table[17] = 36'hF7A385EEF;
        finv_table[16] = 36'hF81F7DEFE;
        finv_table[15] = 36'hF89BB3F0D;
        finv_table[14] = 36'hF91827F1D;
        finv_table[13] = 36'hF994D7F2C;
        finv_table[12] = 36'hFA11C5F3B;
        finv_table[11] = 36'hFA8EF3F4B;
        finv_table[10] = 36'hFB0C5DF5B;
        finv_table[9] = 36'hFB8A05F6A;
        finv_table[8] = 36'hFC07EBF79;
        finv_table[7] = 36'hFC8611F89;
        finv_table[6] = 36'hFD0475F99;
        finv_table[5] = 36'hFD8317FA8;
        finv_table[4] = 36'hFE01F9FB8;
        finv_table[3] = 36'hFE811BFC8;
        finv_table[2] = 36'hFF007BFD8;
        finv_table[1] = 36'hFF801BFE8;
        finv_table[0] = 36'hFFFFFBFF8;
    end

    always @(posedge clk) begin
        dout <= finv_table[addr];
    end

endmodule

`default_nettype wire