module inst_data_mem_blk
(input wire clk,
input wire we,
input wire en,
input wire [31:0] addr,
input wire [31:0] di,
output wire [7:0]
);
