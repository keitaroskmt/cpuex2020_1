`default_nettype none

module fmove
    ( input wire [31:0] x,
      output wire [31:0] y
);
    assign y = x;

endmodule

`default_nettype wire